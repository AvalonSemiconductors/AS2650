magic
tech gf180mcuD
magscale 1 10
timestamp 1701124920
<< metal1 >>
rect 446786 549390 446798 549442
rect 446850 549439 446862 549442
rect 449586 549439 449598 549442
rect 446850 549393 449598 549439
rect 446850 549390 446862 549393
rect 449586 549390 449598 549393
rect 449650 549390 449662 549442
rect 304210 275214 304222 275266
rect 304274 275263 304286 275266
rect 304882 275263 304894 275266
rect 304274 275217 304894 275263
rect 304274 275214 304286 275217
rect 304882 275214 304894 275217
rect 304946 275214 304958 275266
rect 314626 272974 314638 273026
rect 314690 273023 314702 273026
rect 315634 273023 315646 273026
rect 314690 272977 315646 273023
rect 314690 272974 314702 272977
rect 315634 272974 315646 272977
rect 315698 272974 315710 273026
rect 324370 272974 324382 273026
rect 324434 273023 324446 273026
rect 325378 273023 325390 273026
rect 324434 272977 325390 273023
rect 324434 272974 324446 272977
rect 325378 272974 325390 272977
rect 325442 272974 325454 273026
rect 373650 272974 373662 273026
rect 373714 273023 373726 273026
rect 374546 273023 374558 273026
rect 373714 272977 374558 273023
rect 373714 272974 373726 272977
rect 374546 272974 374558 272977
rect 374610 272974 374622 273026
<< via1 >>
rect 446798 549390 446850 549442
rect 449598 549390 449650 549442
rect 304222 275214 304274 275266
rect 304894 275214 304946 275266
rect 314638 272974 314690 273026
rect 315646 272974 315698 273026
rect 324382 272974 324434 273026
rect 325390 272974 325442 273026
rect 373662 272974 373714 273026
rect 374558 272974 374610 273026
<< metal2 >>
rect 11032 595672 11256 597000
rect 11004 595560 11256 595672
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 33096 595560 33348 595672
rect 55160 595560 55412 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 99288 595560 99540 595672
rect 11004 563668 11060 595560
rect 33292 590548 33348 595560
rect 55356 590660 55412 595560
rect 55356 590594 55412 590604
rect 33292 590482 33348 590492
rect 11004 563602 11060 563612
rect 50316 588868 50372 588878
rect 4284 516628 4340 516638
rect 4172 502516 4228 502526
rect 4172 435988 4228 502460
rect 4284 452788 4340 516572
rect 20972 486388 21028 486398
rect 15932 466228 15988 466238
rect 14252 464548 14308 464558
rect 4284 452722 4340 452732
rect 4396 460180 4452 460190
rect 4396 436212 4452 460124
rect 12572 457828 12628 457838
rect 7532 449428 7588 449438
rect 4396 436146 4452 436156
rect 4956 446068 5012 446078
rect 4956 436100 5012 446012
rect 4956 436034 5012 436044
rect 4172 435922 4228 435932
rect 4620 429828 4676 429838
rect 4396 429716 4452 429726
rect 4172 429604 4228 429614
rect 4172 375732 4228 429548
rect 4396 389732 4452 429660
rect 4620 418068 4676 429772
rect 4620 418002 4676 418012
rect 4396 389666 4452 389676
rect 4172 375666 4228 375676
rect 4284 271572 4340 271582
rect 4172 269780 4228 269790
rect 4172 164052 4228 269724
rect 4284 178052 4340 271516
rect 4508 266308 4564 266318
rect 4396 264740 4452 264750
rect 4396 192276 4452 264684
rect 4508 220500 4564 266252
rect 4508 220434 4564 220444
rect 4396 192210 4452 192220
rect 4284 177986 4340 177996
rect 4172 163986 4228 163996
rect 4172 160692 4228 160702
rect 4172 135828 4228 160636
rect 4172 135762 4228 135772
rect 7532 65268 7588 449372
rect 7532 65202 7588 65212
rect 11340 141988 11396 141998
rect 11340 480 11396 141932
rect 12572 93268 12628 457772
rect 12572 93202 12628 93212
rect 14252 50932 14308 464492
rect 14252 50866 14308 50876
rect 15932 8596 15988 466172
rect 19292 446068 19348 446078
rect 15932 8530 15988 8540
rect 17612 211092 17668 211102
rect 15372 4452 15428 4462
rect 13356 4340 13412 4350
rect 13356 480 13412 4284
rect 15372 480 15428 4396
rect 17612 4340 17668 211036
rect 19292 107380 19348 446012
rect 19292 107314 19348 107324
rect 20972 36820 21028 486332
rect 20972 36754 21028 36764
rect 22652 467908 22708 467918
rect 17612 4274 17668 4284
rect 18956 24388 19012 24398
rect 17276 4228 17332 4238
rect 17276 480 17332 4172
rect 11340 392 11592 480
rect 11368 -960 11592 392
rect 13272 -960 13496 480
rect 15176 392 15428 480
rect 17080 392 17332 480
rect 18956 480 19012 24332
rect 22652 22708 22708 467852
rect 50204 420420 50260 420430
rect 48636 416388 48692 416398
rect 48412 401604 48468 401614
rect 26012 286804 26068 286814
rect 22652 22642 22708 22652
rect 24332 231028 24388 231038
rect 20860 13412 20916 13422
rect 20860 480 20916 13356
rect 24332 4228 24388 230972
rect 24332 4162 24388 4172
rect 24668 217700 24724 217710
rect 22988 4116 23044 4126
rect 22988 480 23044 4060
rect 18956 392 19208 480
rect 20860 392 21112 480
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 -960 21112 392
rect 22792 392 23044 480
rect 24668 480 24724 217644
rect 26012 24388 26068 286748
rect 26012 24322 26068 24332
rect 27692 286692 27748 286702
rect 27692 13412 27748 286636
rect 27692 13346 27748 13356
rect 29372 285124 29428 285134
rect 29372 4340 29428 285068
rect 32732 278404 32788 278414
rect 31052 214340 31108 214350
rect 29372 4274 29428 4284
rect 30604 4900 30660 4910
rect 26796 4228 26852 4238
rect 26796 480 26852 4172
rect 30604 480 30660 4844
rect 31052 4116 31108 214284
rect 32732 4900 32788 278348
rect 48412 257908 48468 401548
rect 48412 257842 48468 257852
rect 48524 397572 48580 397582
rect 45612 254548 45668 254558
rect 32732 4834 32788 4844
rect 34412 252868 34468 252878
rect 31052 4050 31108 4060
rect 32508 4340 32564 4350
rect 32508 480 32564 4284
rect 34412 4340 34468 252812
rect 42812 251188 42868 251198
rect 37996 224308 38052 224318
rect 34412 4274 34468 4284
rect 34524 4564 34580 4574
rect 34524 2324 34580 4508
rect 34412 2268 34580 2324
rect 34412 480 34468 2268
rect 37996 480 38052 224252
rect 40124 4900 40180 4910
rect 40124 480 40180 4844
rect 42028 4340 42084 4350
rect 41916 4284 42028 4340
rect 41916 480 41972 4284
rect 42028 4274 42084 4284
rect 42812 4340 42868 251132
rect 44492 232708 44548 232718
rect 44492 4900 44548 232652
rect 44492 4834 44548 4844
rect 42812 4274 42868 4284
rect 45612 480 45668 254492
rect 48524 222740 48580 397516
rect 48524 222674 48580 222684
rect 47852 219268 47908 219278
rect 47852 4340 47908 219212
rect 48636 215908 48692 416332
rect 49980 415044 50036 415054
rect 49980 285012 50036 414988
rect 49980 284946 50036 284956
rect 50092 402948 50148 402958
rect 50092 266420 50148 402892
rect 50092 266354 50148 266364
rect 49532 246148 49588 246158
rect 48636 215842 48692 215852
rect 49420 222628 49476 222638
rect 47852 4274 47908 4284
rect 47740 4228 47796 4238
rect 47740 480 47796 4172
rect 24668 392 24920 480
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 392 26852 480
rect 26600 -960 26824 392
rect 28504 -960 28728 480
rect 30408 392 30660 480
rect 32312 392 32564 480
rect 34216 392 34468 480
rect 30408 -960 30632 392
rect 32312 -960 32536 392
rect 34216 -960 34440 392
rect 36120 -960 36344 480
rect 37996 392 38248 480
rect 38024 -960 38248 392
rect 39928 392 40180 480
rect 39928 -960 40152 392
rect 41832 -960 42056 480
rect 43736 -960 43960 480
rect 45612 392 45864 480
rect 45640 -960 45864 392
rect 47544 392 47796 480
rect 49420 480 49476 222572
rect 49532 4228 49588 246092
rect 50204 227668 50260 420364
rect 50316 342468 50372 588812
rect 55356 583828 55412 583838
rect 53676 582148 53732 582158
rect 51884 578788 51940 578798
rect 50316 342402 50372 342412
rect 51772 398916 51828 398926
rect 51772 283332 51828 398860
rect 51884 314244 51940 578732
rect 51884 314178 51940 314188
rect 51996 432180 52052 432190
rect 51772 283266 51828 283276
rect 50204 227602 50260 227612
rect 51212 234388 51268 234398
rect 51212 4564 51268 234332
rect 51996 160468 52052 432124
rect 53676 339780 53732 582092
rect 53676 339714 53732 339724
rect 55244 430388 55300 430398
rect 53676 324324 53732 324334
rect 51996 160402 52052 160412
rect 53228 229348 53284 229358
rect 51212 4498 51268 4508
rect 49532 4162 49588 4172
rect 53228 480 53284 229292
rect 53676 212660 53732 324268
rect 55244 212884 55300 430332
rect 55356 341124 55412 583772
rect 58716 582260 58772 582270
rect 58492 572180 58548 572190
rect 57036 567028 57092 567038
rect 56924 430164 56980 430174
rect 56812 427364 56868 427374
rect 56700 427252 56756 427262
rect 56700 411012 56756 427196
rect 56700 410946 56756 410956
rect 56812 409668 56868 427308
rect 56812 409602 56868 409612
rect 56924 405636 56980 430108
rect 56924 405570 56980 405580
rect 56924 400260 56980 400270
rect 56700 396228 56756 396238
rect 55356 341058 55412 341068
rect 56252 394884 56308 394894
rect 56252 324324 56308 394828
rect 56700 354452 56756 396172
rect 56700 354386 56756 354396
rect 56812 393540 56868 393550
rect 56252 324258 56308 324268
rect 56812 307412 56868 393484
rect 56812 307346 56868 307356
rect 55244 212818 55300 212828
rect 55356 300804 55412 300814
rect 53676 212594 53732 212604
rect 55356 33684 55412 300748
rect 56700 300804 56756 300814
rect 56700 291844 56756 300748
rect 56924 300132 56980 400204
rect 57036 318276 57092 566972
rect 58380 423108 58436 423118
rect 58268 419076 58324 419086
rect 57036 318210 57092 318220
rect 58156 417732 58212 417742
rect 56924 300066 56980 300076
rect 56700 291778 56756 291788
rect 56812 299460 56868 299470
rect 56812 276500 56868 299404
rect 57036 298116 57092 298126
rect 56812 276434 56868 276444
rect 56924 294084 56980 294094
rect 55356 33618 55412 33628
rect 56252 273140 56308 273150
rect 55356 5012 55412 5022
rect 55356 480 55412 4956
rect 56252 5012 56308 273084
rect 56924 269892 56980 294028
rect 56924 269826 56980 269836
rect 57036 269668 57092 298060
rect 58156 288148 58212 417676
rect 58156 288082 58212 288092
rect 58268 284900 58324 419020
rect 58268 284834 58324 284844
rect 57036 269602 57092 269612
rect 58380 217588 58436 423052
rect 58492 343812 58548 572124
rect 58492 343746 58548 343756
rect 58604 565460 58660 565470
rect 58604 316932 58660 565404
rect 58604 316866 58660 316876
rect 58716 315588 58772 582204
rect 77308 565348 77364 595560
rect 99484 590772 99540 595560
rect 99484 590706 99540 590716
rect 121324 595560 121576 595672
rect 143388 595560 143640 595672
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 165480 595560 165732 595672
rect 121324 570388 121380 595560
rect 121324 570322 121380 570332
rect 121772 572068 121828 572078
rect 77308 565282 77364 565292
rect 104412 488068 104468 488078
rect 101724 437668 101780 437678
rect 99036 434308 99092 434318
rect 90972 432964 91028 432974
rect 66780 432180 66836 432190
rect 64092 432068 64148 432078
rect 60396 431956 60452 431966
rect 60060 425124 60116 425134
rect 58716 315522 58772 315532
rect 59612 354452 59668 354462
rect 58380 217522 58436 217532
rect 58716 286580 58772 286590
rect 58604 214228 58660 214238
rect 56252 4946 56308 4956
rect 57148 139412 57204 139422
rect 57148 480 57204 139356
rect 58604 4004 58660 214172
rect 58716 37940 58772 286524
rect 59612 212772 59668 354396
rect 59836 307412 59892 307422
rect 59612 212706 59668 212716
rect 59724 286468 59780 286478
rect 58716 37874 58772 37884
rect 58940 211204 58996 211214
rect 58604 3938 58660 3948
rect 58940 480 58996 211148
rect 59724 37828 59780 286412
rect 59836 212996 59892 307356
rect 60060 283108 60116 425068
rect 60172 423892 60228 423902
rect 60172 284788 60228 423836
rect 60172 284722 60228 284732
rect 60284 421652 60340 421662
rect 60284 283220 60340 421596
rect 60284 283154 60340 283164
rect 60060 283042 60116 283052
rect 60396 278180 60452 431900
rect 64092 429912 64148 432012
rect 66780 429912 66836 432124
rect 88284 432068 88340 432078
rect 72156 431956 72212 431966
rect 69468 430276 69524 430286
rect 69468 429912 69524 430220
rect 72156 429912 72212 431900
rect 82908 431956 82964 431966
rect 77532 431844 77588 431854
rect 77532 429912 77588 431788
rect 82908 429912 82964 431900
rect 85596 431956 85652 431966
rect 85596 429912 85652 431900
rect 88284 429912 88340 432012
rect 90972 429912 91028 432908
rect 96348 432628 96404 432638
rect 93660 430276 93716 430286
rect 93660 429912 93716 430220
rect 96348 429912 96404 432572
rect 99036 429912 99092 434252
rect 101724 429912 101780 437612
rect 104412 429912 104468 488012
rect 109788 484708 109844 484718
rect 107100 432740 107156 432750
rect 107100 429912 107156 432684
rect 109788 429912 109844 484652
rect 120540 469588 120596 469598
rect 117852 433524 117908 433534
rect 112476 432292 112532 432302
rect 112476 429912 112532 432236
rect 115164 432180 115220 432190
rect 115164 429912 115220 432124
rect 117852 429912 117908 433468
rect 120540 429912 120596 469532
rect 121772 432740 121828 572012
rect 143388 555268 143444 595560
rect 165676 590884 165732 595560
rect 165676 590818 165732 590828
rect 187516 595560 187768 595672
rect 209608 595672 209832 597000
rect 209608 595560 209860 595672
rect 231672 595560 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 253736 595560 253988 595672
rect 275800 595560 276052 595672
rect 297864 595560 298116 595672
rect 319928 595560 320180 595672
rect 143388 555202 143444 555212
rect 153692 557844 153748 557854
rect 144732 500724 144788 500734
rect 136668 499828 136724 499838
rect 133980 498148 134036 498158
rect 131292 437780 131348 437790
rect 121772 432674 121828 432684
rect 123228 433636 123284 433646
rect 123228 429912 123284 433580
rect 128604 432404 128660 432414
rect 128604 429912 128660 432348
rect 131292 429912 131348 437724
rect 133980 429912 134036 498092
rect 136668 429912 136724 499772
rect 142044 434532 142100 434542
rect 139356 434420 139412 434430
rect 139356 429912 139412 434364
rect 142044 429912 142100 434476
rect 144732 429912 144788 500668
rect 150108 498260 150164 498270
rect 147420 494788 147476 494798
rect 147420 429912 147476 494732
rect 150108 429912 150164 498204
rect 153692 476308 153748 557788
rect 173740 557844 173796 557854
rect 173740 554904 173796 557788
rect 187516 555380 187572 595560
rect 209804 590996 209860 595560
rect 231756 591108 231812 595560
rect 231756 591042 231812 591052
rect 209804 590930 209860 590940
rect 253932 588980 253988 595560
rect 275996 590212 276052 595560
rect 298060 591220 298116 595560
rect 320124 591332 320180 595560
rect 320124 591266 320180 591276
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 430220 595560 430472 595672
rect 452284 595560 452536 595672
rect 474348 595560 474600 595672
rect 496412 595560 496664 595672
rect 518476 595560 518728 595672
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 298060 591154 298116 591164
rect 279692 590996 279748 591006
rect 275996 590146 276052 590156
rect 278012 590212 278068 590222
rect 253932 588914 253988 588924
rect 187516 555314 187572 555324
rect 274652 554484 274708 554494
rect 201292 554372 201348 554382
rect 201292 554306 201348 554316
rect 216748 551572 216804 551582
rect 215740 548884 215796 548894
rect 215180 543508 215236 543518
rect 214508 510804 214564 510814
rect 214396 505764 214452 505774
rect 160860 501508 160916 501518
rect 153692 476242 153748 476252
rect 155484 499940 155540 499950
rect 152796 444388 152852 444398
rect 152796 429912 152852 444332
rect 155484 429912 155540 499884
rect 158172 437892 158228 437902
rect 158172 429912 158228 437836
rect 160860 429912 160916 501452
rect 176988 500612 177044 500622
rect 162764 486388 162820 500136
rect 162764 486322 162820 486332
rect 167244 446068 167300 500136
rect 167244 446002 167300 446012
rect 171500 500052 171556 500062
rect 163548 433412 163604 433422
rect 163548 429912 163604 433356
rect 166236 433412 166292 433422
rect 166236 429912 166292 433356
rect 169596 433412 169652 433422
rect 169596 429940 169652 433356
rect 168952 429884 169652 429940
rect 171500 429940 171556 499996
rect 171724 449428 171780 500136
rect 176204 467908 176260 500136
rect 176204 467842 176260 467852
rect 171724 449362 171780 449372
rect 174300 449428 174356 449438
rect 171500 429884 171640 429940
rect 174300 429912 174356 449372
rect 176988 429912 177044 500556
rect 179676 493108 179732 493118
rect 179676 429912 179732 493052
rect 180684 457828 180740 500136
rect 180684 457762 180740 457772
rect 182364 491428 182420 491438
rect 182364 429912 182420 491372
rect 185164 464548 185220 500136
rect 189644 466228 189700 500136
rect 194124 496468 194180 500136
rect 198604 496580 198660 500136
rect 198604 496514 198660 496524
rect 202412 500108 203112 500164
rect 202412 497252 202468 500108
rect 194124 496402 194180 496412
rect 189644 466162 189700 466172
rect 185164 464482 185220 464492
rect 187740 451108 187796 451118
rect 185052 438004 185108 438014
rect 185052 429912 185108 437948
rect 187740 429912 187796 451052
rect 202412 444388 202468 497196
rect 207564 452900 207620 500136
rect 212044 469588 212100 500136
rect 212044 469522 212100 469532
rect 207564 452834 207620 452844
rect 202412 444322 202468 444332
rect 190428 439348 190484 439358
rect 190428 429912 190484 439292
rect 214396 437892 214452 505708
rect 214396 437826 214452 437836
rect 214508 437780 214564 510748
rect 215068 508564 215124 508574
rect 214844 502852 214900 502862
rect 214844 499940 214900 502796
rect 215068 501508 215124 508508
rect 215068 501442 215124 501452
rect 214844 499874 214900 499884
rect 215180 491428 215236 543452
rect 215292 540820 215348 540830
rect 215292 493108 215348 540764
rect 215404 538132 215460 538142
rect 215404 501732 215460 538076
rect 215404 501666 215460 501676
rect 215516 516628 215572 516638
rect 215516 499828 215572 516572
rect 215516 499762 215572 499772
rect 215628 513940 215684 513950
rect 215628 513268 215684 513884
rect 215628 498148 215684 513212
rect 215628 498082 215684 498092
rect 215292 493042 215348 493052
rect 215180 491362 215236 491372
rect 215740 451108 215796 548828
rect 215740 451042 215796 451052
rect 216748 439348 216804 551516
rect 217532 550228 217588 550238
rect 217308 532756 217364 532766
rect 217084 530068 217140 530078
rect 216748 439282 216804 439292
rect 216860 521668 216916 521678
rect 214508 437714 214564 437724
rect 216860 434532 216916 521612
rect 216860 434466 216916 434476
rect 216972 519988 217028 519998
rect 216972 434420 217028 519932
rect 217084 498260 217140 530012
rect 217084 498194 217140 498204
rect 217196 527492 217252 527502
rect 217196 494788 217252 527436
rect 217308 501620 217364 532700
rect 217308 501554 217364 501564
rect 217532 524692 217588 550172
rect 217756 549444 217812 549454
rect 217756 527492 217812 549388
rect 217756 527426 217812 527436
rect 218428 546196 218484 546206
rect 217532 500724 217588 524636
rect 217532 500658 217588 500668
rect 217196 494722 217252 494732
rect 218428 438004 218484 546140
rect 218540 535444 218596 535454
rect 218540 449428 218596 535388
rect 218540 449362 218596 449372
rect 246876 452900 246932 452910
rect 218428 437938 218484 437948
rect 216972 434354 217028 434364
rect 209244 432628 209300 432638
rect 206556 432516 206612 432526
rect 203868 430612 203924 430622
rect 193116 430388 193172 430398
rect 193116 429912 193172 430332
rect 201180 430388 201236 430398
rect 201180 429912 201236 430332
rect 203868 429912 203924 430556
rect 206556 429912 206612 432460
rect 209244 429912 209300 432572
rect 244188 430836 244244 430846
rect 219996 430724 220052 430734
rect 214620 430500 214676 430510
rect 212828 430052 212884 430062
rect 212716 429996 212828 430052
rect 212716 429940 212772 429996
rect 212828 429986 212884 429996
rect 211960 429884 212772 429940
rect 214620 429912 214676 430444
rect 219996 429912 220052 430668
rect 244188 429912 244244 430780
rect 246876 429912 246932 452844
rect 265692 433412 265748 433422
rect 257628 431060 257684 431070
rect 254940 430948 254996 430958
rect 254940 429912 254996 430892
rect 257628 429912 257684 431004
rect 265692 429912 265748 433356
rect 268716 433412 268772 433422
rect 268716 429940 268772 433356
rect 268408 429884 268772 429940
rect 272636 432740 272692 432750
rect 80220 429492 80276 429502
rect 80220 429426 80276 429436
rect 74844 429380 74900 429390
rect 74844 429314 74900 429324
rect 125916 429268 125972 429278
rect 60620 429212 61432 429268
rect 60620 428596 60676 429212
rect 125916 429202 125972 429212
rect 217308 429268 217364 429278
rect 217308 429202 217364 429212
rect 249564 429268 249620 429278
rect 249564 429202 249620 429212
rect 252252 429268 252308 429278
rect 252252 429202 252308 429212
rect 260316 429268 260372 429278
rect 260316 429202 260372 429212
rect 263004 429268 263060 429278
rect 263004 429202 263060 429212
rect 60620 428530 60676 428540
rect 270620 422436 270676 422446
rect 269500 410004 269556 410014
rect 269388 405748 269444 405758
rect 60396 278114 60452 278124
rect 60620 300132 60676 300142
rect 59836 212930 59892 212940
rect 60620 212548 60676 300076
rect 63756 290164 63812 290174
rect 62972 290108 63756 290164
rect 60620 212482 60676 212492
rect 61180 286916 61236 286926
rect 60284 210980 60340 210990
rect 60172 210868 60228 210878
rect 59724 37762 59780 37772
rect 59948 209524 60004 209534
rect 59948 4340 60004 209468
rect 59948 4274 60004 4284
rect 60060 209412 60116 209422
rect 60060 4116 60116 209356
rect 60172 4452 60228 210812
rect 60172 4386 60228 4396
rect 60284 4228 60340 210924
rect 61180 139412 61236 286860
rect 62972 209972 63028 290108
rect 63756 290098 63812 290108
rect 65212 211092 65268 290136
rect 67228 285124 67284 290136
rect 67228 285058 67284 285068
rect 69244 231028 69300 290136
rect 71260 286804 71316 290136
rect 71260 286738 71316 286748
rect 73276 286692 73332 290136
rect 73276 286626 73332 286636
rect 69244 230962 69300 230972
rect 75292 214340 75348 290136
rect 77308 217700 77364 290136
rect 79324 219268 79380 290136
rect 81340 278404 81396 290136
rect 81340 278338 81396 278348
rect 83356 252868 83412 290136
rect 83356 252802 83412 252812
rect 85372 234388 85428 290136
rect 85372 234322 85428 234332
rect 87388 224308 87444 290136
rect 89404 232708 89460 290136
rect 89404 232642 89460 232652
rect 91196 283332 91252 283342
rect 87388 224242 87444 224252
rect 79324 219202 79380 219212
rect 87164 222740 87220 222750
rect 77308 217634 77364 217644
rect 75292 214274 75348 214284
rect 65212 211026 65268 211036
rect 66668 213332 66724 213342
rect 66668 209972 66724 213276
rect 75068 212996 75124 213006
rect 71036 212884 71092 212894
rect 66668 209916 67032 209972
rect 71036 209944 71092 212828
rect 75068 209944 75124 212940
rect 83132 212772 83188 212782
rect 79100 212660 79156 212670
rect 79100 209944 79156 212604
rect 83132 209944 83188 212716
rect 87164 209944 87220 222684
rect 91196 209944 91252 283276
rect 91420 251188 91476 290136
rect 93436 254548 93492 290136
rect 93436 254482 93492 254492
rect 91420 251122 91476 251132
rect 95452 246148 95508 290136
rect 95452 246082 95508 246092
rect 96572 285684 96628 285694
rect 96572 222628 96628 285628
rect 97468 285684 97524 290136
rect 97468 285618 97524 285628
rect 96572 222562 96628 222572
rect 99260 257908 99316 257918
rect 95228 212548 95284 212558
rect 95228 209944 95284 212492
rect 99260 209944 99316 257852
rect 99484 229348 99540 290136
rect 101500 273140 101556 290136
rect 103516 286916 103572 290136
rect 103516 286850 103572 286860
rect 101500 273074 101556 273084
rect 99484 229282 99540 229292
rect 103292 266420 103348 266430
rect 103292 209944 103348 266364
rect 105532 211204 105588 290136
rect 105532 211138 105588 211148
rect 107324 285012 107380 285022
rect 107324 209944 107380 284956
rect 62972 209906 63028 209916
rect 107548 209524 107604 290136
rect 107548 209458 107604 209468
rect 109564 209412 109620 290136
rect 111356 215908 111412 215918
rect 111356 209944 111412 215852
rect 111580 210980 111636 290136
rect 111580 210914 111636 210924
rect 113596 210868 113652 290136
rect 113596 210802 113652 210812
rect 115388 288148 115444 288158
rect 115388 209944 115444 288092
rect 115612 281428 115668 290136
rect 115612 281362 115668 281372
rect 117628 227780 117684 290136
rect 119644 286580 119700 290136
rect 119644 286514 119700 286524
rect 117628 227714 117684 227724
rect 119420 284900 119476 284910
rect 119420 209944 119476 284844
rect 121660 214228 121716 290136
rect 123676 286468 123732 290136
rect 123676 286402 123732 286412
rect 125692 285684 125748 290136
rect 127708 286356 127764 290136
rect 127708 286290 127764 286300
rect 125692 285618 125748 285628
rect 127484 283220 127540 283230
rect 121660 214162 121716 214172
rect 123452 227668 123508 227678
rect 123452 209944 123508 227612
rect 127484 209944 127540 283164
rect 129724 258020 129780 290136
rect 131740 286580 131796 290136
rect 131740 286514 131796 286524
rect 129724 257954 129780 257964
rect 133756 231140 133812 290136
rect 135772 286356 135828 290136
rect 135772 286290 135828 286300
rect 137788 286244 137844 290136
rect 137788 286178 137844 286188
rect 139804 285684 139860 290136
rect 139804 285618 139860 285628
rect 141820 285684 141876 290136
rect 143836 286580 143892 290136
rect 143836 286514 143892 286524
rect 145852 286020 145908 290136
rect 147868 286244 147924 290136
rect 147868 286178 147924 286188
rect 145852 285954 145908 285964
rect 149884 285796 149940 290136
rect 149884 285730 149940 285740
rect 141820 285618 141876 285628
rect 151900 285124 151956 290136
rect 153916 285684 153972 290136
rect 153916 285618 153972 285628
rect 155932 285684 155988 290136
rect 155932 285618 155988 285628
rect 157052 285684 157108 285694
rect 151900 285058 151956 285068
rect 151676 284900 151732 284910
rect 133756 231074 133812 231084
rect 135548 284788 135604 284798
rect 131516 217588 131572 217598
rect 131516 209944 131572 217532
rect 135548 209944 135604 284732
rect 143612 284788 143668 284798
rect 139580 283108 139636 283118
rect 139580 209944 139636 283052
rect 143612 209944 143668 284732
rect 147644 283108 147700 283118
rect 147644 209944 147700 283052
rect 151676 209944 151732 284844
rect 157052 222628 157108 285628
rect 157948 285684 158004 290136
rect 157948 285618 158004 285628
rect 159740 290108 159992 290164
rect 159740 285684 159796 290108
rect 159740 285618 159796 285628
rect 157052 222562 157108 222572
rect 155708 217588 155764 217598
rect 155708 209944 155764 217532
rect 159740 212548 159796 212558
rect 159740 209944 159796 212492
rect 109564 209346 109620 209356
rect 161980 209412 162036 290136
rect 163996 283332 164052 290136
rect 166012 285684 166068 290136
rect 166012 285618 166068 285628
rect 163996 283266 164052 283276
rect 167804 266420 167860 266430
rect 163772 222628 163828 222638
rect 163772 209944 163828 222572
rect 167804 209944 167860 266364
rect 168028 210868 168084 290136
rect 170044 286916 170100 290136
rect 170044 286850 170100 286860
rect 172060 212772 172116 290136
rect 174076 285684 174132 290136
rect 174076 285618 174132 285628
rect 176092 285684 176148 290136
rect 176092 285618 176148 285628
rect 178108 285684 178164 290136
rect 178108 285618 178164 285628
rect 180124 231028 180180 290136
rect 180124 230962 180180 230972
rect 179900 212884 179956 212894
rect 172060 212706 172116 212716
rect 175868 212772 175924 212782
rect 168028 210802 168084 210812
rect 171836 212660 171892 212670
rect 171836 209944 171892 212604
rect 175868 209944 175924 212716
rect 179900 209944 179956 212828
rect 182140 210980 182196 290136
rect 184156 285684 184212 290136
rect 184156 285618 184212 285628
rect 186172 285684 186228 290136
rect 186172 285618 186228 285628
rect 188188 285684 188244 290136
rect 190204 286468 190260 290136
rect 190204 286402 190260 286412
rect 191548 290108 192248 290164
rect 188188 285618 188244 285628
rect 191548 285684 191604 290108
rect 194236 286692 194292 290136
rect 194236 286626 194292 286636
rect 191548 285618 191604 285628
rect 196252 285684 196308 290136
rect 196252 285618 196308 285628
rect 198268 285684 198324 290136
rect 200284 287028 200340 290136
rect 200284 286962 200340 286972
rect 202300 285796 202356 290136
rect 202300 285730 202356 285740
rect 198268 285618 198324 285628
rect 204316 285684 204372 290136
rect 206332 286804 206388 290136
rect 206332 286738 206388 286748
rect 204316 285618 204372 285628
rect 208348 285684 208404 290136
rect 210364 286916 210420 290136
rect 210364 286850 210420 286860
rect 212380 286580 212436 290136
rect 212380 286514 212436 286524
rect 208348 285618 208404 285628
rect 214396 285684 214452 290136
rect 214396 285618 214452 285628
rect 216412 285684 216468 290136
rect 216412 285618 216468 285628
rect 218428 285684 218484 290136
rect 220444 286468 220500 290136
rect 220444 286402 220500 286412
rect 221788 290108 222488 290164
rect 218428 285618 218484 285628
rect 221788 285684 221844 290108
rect 221788 285618 221844 285628
rect 196028 285012 196084 285022
rect 191996 283220 192052 283230
rect 187964 224308 188020 224318
rect 182140 210914 182196 210924
rect 183932 214228 183988 214238
rect 183932 209944 183988 214172
rect 187964 209944 188020 224252
rect 191996 209944 192052 283164
rect 196028 209944 196084 284956
rect 200060 283332 200116 283342
rect 200060 209944 200116 283276
rect 224476 281428 224532 290136
rect 226492 285684 226548 290136
rect 226492 285618 226548 285628
rect 228508 285684 228564 290136
rect 230524 285796 230580 290136
rect 230524 285730 230580 285740
rect 231868 290108 232568 290164
rect 228508 285618 228564 285628
rect 231868 285684 231924 290108
rect 231868 285618 231924 285628
rect 224476 281362 224532 281372
rect 228284 261380 228340 261390
rect 222572 260484 222628 260494
rect 216188 259700 216244 259710
rect 208124 258804 208180 258814
rect 204092 257908 204148 257918
rect 204092 209944 204148 257852
rect 208124 209944 208180 258748
rect 212156 215908 212212 215918
rect 212156 209944 212212 215852
rect 216188 209944 216244 259644
rect 220220 213332 220276 213342
rect 220220 209944 220276 213276
rect 222572 213332 222628 260428
rect 222572 213266 222628 213276
rect 224252 259812 224308 259822
rect 224252 209944 224308 259756
rect 228284 209944 228340 261324
rect 232316 258916 232372 258926
rect 232316 209944 232372 258860
rect 234556 210868 234612 290136
rect 236572 286468 236628 290136
rect 236572 286402 236628 286412
rect 238588 285684 238644 290136
rect 238588 285618 238644 285628
rect 240604 285684 240660 290136
rect 240604 285618 240660 285628
rect 242620 285684 242676 290136
rect 244636 285796 244692 290136
rect 246680 290108 246932 290164
rect 248696 290108 249284 290164
rect 244636 285730 244692 285740
rect 242620 285618 242676 285628
rect 246876 285684 246932 290108
rect 246876 285618 246932 285628
rect 249228 285684 249284 290108
rect 250684 286356 250740 290136
rect 250684 286290 250740 286300
rect 252140 290108 252728 290164
rect 249228 285618 249284 285628
rect 252140 285684 252196 290108
rect 254716 286468 254772 290136
rect 254716 286402 254772 286412
rect 252140 285618 252196 285628
rect 256732 285684 256788 290136
rect 256732 285618 256788 285628
rect 258748 285684 258804 290136
rect 258748 285618 258804 285628
rect 260428 290108 260792 290164
rect 260428 285684 260484 290108
rect 262780 285908 262836 290136
rect 262780 285842 262836 285852
rect 264796 285796 264852 290136
rect 264796 285730 264852 285740
rect 260428 285618 260484 285628
rect 266812 285684 266868 290136
rect 266812 285618 266868 285628
rect 248444 270004 248500 270014
rect 234556 210802 234612 210812
rect 236348 261492 236404 261502
rect 236348 209944 236404 261436
rect 240380 254548 240436 254558
rect 240380 209944 240436 254492
rect 244412 217700 244468 217710
rect 244412 209944 244468 217644
rect 248444 209944 248500 269948
rect 264572 268212 264628 268222
rect 260540 222740 260596 222750
rect 256508 216020 256564 216030
rect 252476 214340 252532 214350
rect 252476 209944 252532 214284
rect 256508 209944 256564 215964
rect 260540 209944 260596 222684
rect 264572 209944 264628 268156
rect 268604 266532 268660 266542
rect 268604 209944 268660 266476
rect 269388 217588 269444 405692
rect 269500 266420 269556 409948
rect 270508 408996 270564 409006
rect 269500 266354 269556 266364
rect 269612 347844 269668 347854
rect 269388 217522 269444 217532
rect 269612 212548 269668 347788
rect 269836 306292 269892 306302
rect 269724 304052 269780 304062
rect 269724 289828 269780 303996
rect 269724 289762 269780 289772
rect 269836 212772 269892 306236
rect 270508 222628 270564 408940
rect 270620 257908 270676 422380
rect 270732 421092 270788 421102
rect 270732 283332 270788 421036
rect 270844 419748 270900 419758
rect 270844 285012 270900 419692
rect 272188 414372 272244 414382
rect 270844 284946 270900 284956
rect 270956 404964 271012 404974
rect 270956 284900 271012 404908
rect 270956 284834 271012 284844
rect 271292 334404 271348 334414
rect 270732 283266 270788 283276
rect 270620 257842 270676 257852
rect 270508 222562 270564 222572
rect 269836 212706 269892 212716
rect 271292 212660 271348 334348
rect 272188 302428 272244 414316
rect 272300 413028 272356 413038
rect 272300 306292 272356 412972
rect 272412 411684 272468 411694
rect 272412 334404 272468 411628
rect 272524 407652 272580 407662
rect 272524 347844 272580 407596
rect 272636 388836 272692 432684
rect 272972 432628 273028 432638
rect 272972 397348 273028 432572
rect 273980 418404 274036 418414
rect 272972 397282 273028 397292
rect 273868 415716 273924 415726
rect 272636 388770 272692 388780
rect 272972 381444 273028 381454
rect 272972 370020 273028 381388
rect 272972 369954 273028 369964
rect 272524 347778 272580 347788
rect 272412 334338 272468 334348
rect 273084 335076 273140 335086
rect 272300 306226 272356 306236
rect 272972 333732 273028 333742
rect 271516 302372 272244 302428
rect 272300 302820 272356 302830
rect 271516 212884 271572 302372
rect 272300 291508 272356 302764
rect 272300 291442 272356 291452
rect 272972 257908 273028 333676
rect 273084 279748 273140 335020
rect 273084 279682 273140 279692
rect 273196 332388 273252 332398
rect 273196 276612 273252 332332
rect 273196 276546 273252 276556
rect 273308 328356 273364 328366
rect 273308 273252 273364 328300
rect 273532 327012 273588 327022
rect 273420 325668 273476 325678
rect 273420 278404 273476 325612
rect 273532 279860 273588 326956
rect 273756 318948 273812 318958
rect 273756 279972 273812 318892
rect 273756 279906 273812 279916
rect 273532 279794 273588 279804
rect 273420 278338 273476 278348
rect 273308 273186 273364 273196
rect 272972 257842 273028 257852
rect 273868 214228 273924 415660
rect 273980 283220 274036 418348
rect 274092 402276 274148 402286
rect 274092 284788 274148 402220
rect 274652 398244 274708 554428
rect 274652 398178 274708 398188
rect 274764 432516 274820 432526
rect 274764 383908 274820 432460
rect 274764 383842 274820 383852
rect 275548 417060 275604 417070
rect 274092 284722 274148 284732
rect 273980 283154 274036 283164
rect 275548 224308 275604 417004
rect 275660 403620 275716 403630
rect 275660 283108 275716 403564
rect 278012 380212 278068 590156
rect 278124 553588 278180 553598
rect 278124 400932 278180 553532
rect 278124 400866 278180 400876
rect 279692 381892 279748 590940
rect 299964 590996 300020 591006
rect 298284 590436 298340 590446
rect 279804 562212 279860 562222
rect 279804 434308 279860 562156
rect 291452 553476 291508 553486
rect 289772 552916 289828 552926
rect 279804 434242 279860 434252
rect 284732 496580 284788 496590
rect 279692 381826 279748 381836
rect 279804 431956 279860 431966
rect 279804 380548 279860 431900
rect 284732 402948 284788 496524
rect 288092 496468 288148 496478
rect 284732 402882 284788 402892
rect 284844 432292 284900 432302
rect 279804 380482 279860 380492
rect 278012 380146 278068 380156
rect 284844 379652 284900 432236
rect 288092 402836 288148 496412
rect 288092 402770 288148 402780
rect 289772 390180 289828 552860
rect 291452 399588 291508 553420
rect 296492 549780 296548 549790
rect 291452 399522 291508 399532
rect 293132 549668 293188 549678
rect 293132 396900 293188 549612
rect 293132 396834 293188 396844
rect 294812 549332 294868 549342
rect 294812 394212 294868 549276
rect 294812 394146 294868 394156
rect 294924 474292 294980 474302
rect 289772 390114 289828 390124
rect 284844 379586 284900 379596
rect 294924 379540 294980 474236
rect 295036 433636 295092 433646
rect 295036 398132 295092 433580
rect 295260 433524 295316 433534
rect 295148 432180 295204 432190
rect 295148 401492 295204 432124
rect 295148 401426 295204 401436
rect 295260 399812 295316 433468
rect 295260 399746 295316 399756
rect 295036 398066 295092 398076
rect 296492 392868 296548 549724
rect 298172 548772 298228 548782
rect 298060 429828 298116 429838
rect 298060 401380 298116 429772
rect 298060 401314 298116 401324
rect 296492 392802 296548 392812
rect 298172 391524 298228 548716
rect 298284 484708 298340 590380
rect 299852 551124 299908 551134
rect 298284 484642 298340 484652
rect 298396 488404 298452 488414
rect 298172 391458 298228 391468
rect 298284 432404 298340 432414
rect 298284 380100 298340 432348
rect 298396 401268 298452 488348
rect 298844 436100 298900 436110
rect 298620 435988 298676 435998
rect 298396 401202 298452 401212
rect 298508 429716 298564 429726
rect 298508 380324 298564 429660
rect 298620 402612 298676 435932
rect 298620 402546 298676 402556
rect 298844 402276 298900 436044
rect 298844 402210 298900 402220
rect 299852 395556 299908 551068
rect 299964 488068 300020 590940
rect 341964 572180 342020 595560
rect 341964 572114 342020 572124
rect 364028 567028 364084 595560
rect 386092 590436 386148 595560
rect 386092 590370 386148 590380
rect 408268 588868 408324 595560
rect 408268 588802 408324 588812
rect 364028 566962 364084 566972
rect 430220 565460 430276 595560
rect 451276 591220 451332 591230
rect 430220 565394 430276 565404
rect 449372 591108 449428 591118
rect 416780 554484 416836 554494
rect 318220 553364 318276 553374
rect 313292 553252 313348 553262
rect 303436 553140 303492 553150
rect 303436 549864 303492 553084
rect 308364 553028 308420 553038
rect 308364 549864 308420 552972
rect 313292 549864 313348 553196
rect 318220 549864 318276 553308
rect 382396 551572 382452 551582
rect 377356 551460 377412 551470
rect 372428 551348 372484 551358
rect 367500 551236 367556 551246
rect 367164 550004 367220 550014
rect 367164 549892 367220 549948
rect 367500 549892 367556 551180
rect 367164 549864 367556 549892
rect 372428 549892 372484 551292
rect 367164 549836 367528 549864
rect 377356 550228 377412 551404
rect 377356 549864 377412 550172
rect 372428 549826 372484 549836
rect 362572 549556 362628 549566
rect 362572 549490 362628 549500
rect 323148 549444 323204 549454
rect 323148 549378 323204 549388
rect 328076 549444 328132 549454
rect 328076 549378 328132 549388
rect 333004 549444 333060 549454
rect 333004 549378 333060 549388
rect 337932 549444 337988 549454
rect 337932 549378 337988 549388
rect 342860 549444 342916 549454
rect 342860 549378 342916 549388
rect 347788 549444 347844 549454
rect 347788 549378 347844 549388
rect 352716 549444 352772 549454
rect 352716 549378 352772 549388
rect 357644 549444 357700 549454
rect 357644 549378 357700 549388
rect 382284 549444 382340 549454
rect 382396 549444 382452 551516
rect 406924 551124 406980 551134
rect 397068 549892 397124 549902
rect 406924 549864 406980 551068
rect 416780 549864 416836 554428
rect 426636 553588 426692 553598
rect 421708 553476 421764 553486
rect 421708 549864 421764 553420
rect 426636 549864 426692 553532
rect 436492 552916 436548 552926
rect 430780 550116 430836 550126
rect 430780 549892 430836 550060
rect 430780 549836 431592 549892
rect 436492 549864 436548 552860
rect 397068 549826 397124 549836
rect 387212 549780 387268 549790
rect 387212 549714 387268 549724
rect 392812 549780 392868 549790
rect 382340 549388 382452 549444
rect 392140 549444 392196 549454
rect 382284 549378 382340 549388
rect 392140 549378 392196 549388
rect 392812 549444 392868 549724
rect 411852 549668 411908 549678
rect 411852 549602 411908 549612
rect 392812 549378 392868 549388
rect 401996 549332 402052 549342
rect 401996 549266 402052 549276
rect 431340 549332 431396 549836
rect 446796 549444 446852 549454
rect 446376 549442 446852 549444
rect 446376 549390 446798 549442
rect 446850 549390 446852 549442
rect 446376 549388 446852 549390
rect 446796 549378 446852 549388
rect 431340 549266 431396 549276
rect 441420 549332 441476 549342
rect 441420 549266 441476 549276
rect 301084 549108 301140 549118
rect 300972 548660 301028 548670
rect 300972 530068 301028 548604
rect 300972 530002 301028 530012
rect 301084 508228 301140 549052
rect 301084 508162 301140 508172
rect 299964 488002 300020 488012
rect 449372 434420 449428 591052
rect 451052 590548 451108 590558
rect 449372 434354 449428 434364
rect 449484 553140 449540 553150
rect 301084 430836 301140 430846
rect 300860 427700 300916 427710
rect 300860 401156 300916 427644
rect 300860 401090 300916 401100
rect 301084 400484 301140 430780
rect 449484 429604 449540 553084
rect 449596 549442 449652 549454
rect 449596 549390 449598 549442
rect 449650 549390 449652 549442
rect 449596 549388 449652 549390
rect 449596 549332 449764 549388
rect 449708 449428 449764 549332
rect 449708 449362 449764 449372
rect 451052 446180 451108 590492
rect 451052 446114 451108 446124
rect 451164 553252 451220 553262
rect 451164 437668 451220 553196
rect 451276 449540 451332 591164
rect 452284 572068 452340 595560
rect 464492 591332 464548 591342
rect 456204 590884 456260 590894
rect 456092 587188 456148 587198
rect 452284 572002 452340 572012
rect 452732 573076 452788 573086
rect 451276 449474 451332 449484
rect 451164 437602 451220 437612
rect 452732 434308 452788 573020
rect 454412 563668 454468 563678
rect 452844 553364 452900 553374
rect 452844 446068 452900 553308
rect 452844 446002 452900 446012
rect 452732 434242 452788 434252
rect 449484 429538 449540 429548
rect 301084 400418 301140 400428
rect 299852 395490 299908 395500
rect 298508 380258 298564 380268
rect 298284 380034 298340 380044
rect 294924 379474 294980 379484
rect 299068 378980 299124 378990
rect 299068 376740 299124 378924
rect 454412 377636 454468 563612
rect 454524 553028 454580 553038
rect 454524 439348 454580 552972
rect 454524 439282 454580 439292
rect 456092 437892 456148 587132
rect 456204 444388 456260 590828
rect 456204 444322 456260 444332
rect 457772 590772 457828 590782
rect 456092 437826 456148 437836
rect 457772 437780 457828 590716
rect 459564 590660 459620 590670
rect 459452 549332 459508 549342
rect 459452 448532 459508 549276
rect 459564 449652 459620 590604
rect 462812 588980 462868 588990
rect 461244 570388 461300 570398
rect 459564 449586 459620 449596
rect 461132 565348 461188 565358
rect 459452 448466 459508 448476
rect 457772 437714 457828 437724
rect 454412 377570 454468 377580
rect 456092 430052 456148 430062
rect 299068 376674 299124 376684
rect 294924 375396 294980 375406
rect 289772 374052 289828 374062
rect 284732 331044 284788 331054
rect 279020 309540 279076 309550
rect 278908 306852 278964 306862
rect 278796 305508 278852 305518
rect 275660 283042 275716 283052
rect 277676 300132 277732 300142
rect 275548 224242 275604 224252
rect 276668 264964 276724 264974
rect 273868 214162 273924 214172
rect 271516 212818 271572 212828
rect 271292 212594 271348 212604
rect 269612 212482 269668 212492
rect 272636 212548 272692 212558
rect 272636 209944 272692 212492
rect 276668 209944 276724 264908
rect 161980 209346 162036 209356
rect 63672 160076 63812 160132
rect 63756 156324 63812 160076
rect 66332 156548 66388 160104
rect 69020 157780 69076 160104
rect 69020 157714 69076 157724
rect 71708 157108 71764 160104
rect 71708 157042 71764 157052
rect 73836 157780 73892 157790
rect 66332 156482 66388 156492
rect 70476 156548 70532 156558
rect 63756 156268 63924 156324
rect 63868 155540 63924 156268
rect 63868 155474 63924 155484
rect 70476 152180 70532 156492
rect 73836 155428 73892 157724
rect 74396 157220 74452 160104
rect 74396 157154 74452 157164
rect 73836 155362 73892 155372
rect 70476 152114 70532 152124
rect 65436 150388 65492 150398
rect 64428 142324 64484 142334
rect 61180 139346 61236 139356
rect 63756 141204 63812 141214
rect 63756 139048 63812 141148
rect 64428 139048 64484 142268
rect 65436 139076 65492 150332
rect 77084 148708 77140 160104
rect 77084 148642 77140 148652
rect 76076 147028 76132 147038
rect 65352 139020 65492 139076
rect 73500 145460 73556 145470
rect 73500 139048 73556 145404
rect 74620 142212 74676 142222
rect 74172 141988 74228 141998
rect 74172 139048 74228 141932
rect 74620 139048 74676 142156
rect 75068 142100 75124 142110
rect 75068 139048 75124 142044
rect 75516 141316 75572 141326
rect 75516 139048 75572 141260
rect 76076 139048 76132 146972
rect 79772 142100 79828 160104
rect 82460 142212 82516 160104
rect 84924 160076 85176 160132
rect 82460 142146 82516 142156
rect 84252 143668 84308 143678
rect 79772 142034 79828 142044
rect 84252 139048 84308 143612
rect 84924 142324 84980 160076
rect 84924 142258 84980 142268
rect 85036 148708 85092 148718
rect 85036 141092 85092 148652
rect 87836 143780 87892 160104
rect 90524 145572 90580 160104
rect 93212 155764 93268 160104
rect 93212 155698 93268 155708
rect 90524 145506 90580 145516
rect 87836 143714 87892 143724
rect 90972 141764 91028 141774
rect 85036 139048 85092 141036
rect 85820 141428 85876 141438
rect 85820 139048 85876 141372
rect 90972 139048 91028 141708
rect 95900 141764 95956 160104
rect 96908 155540 96964 155550
rect 95900 141698 95956 141708
rect 96460 141764 96516 141774
rect 91980 141540 92036 141550
rect 91980 139048 92036 141484
rect 92764 141204 92820 141214
rect 92764 139048 92820 141148
rect 93324 140644 93380 140654
rect 93324 139048 93380 140588
rect 96460 140308 96516 141708
rect 96460 140242 96516 140252
rect 96908 139300 96964 155484
rect 97692 141540 97748 141550
rect 97692 140420 97748 141484
rect 98588 141540 98644 160104
rect 98588 141474 98644 141484
rect 100828 160076 101304 160132
rect 100828 141204 100884 160076
rect 100828 140532 100884 141148
rect 103964 140644 104020 160104
rect 106680 160076 106820 160132
rect 103964 140578 104020 140588
rect 106652 155652 106708 155662
rect 100828 140466 100884 140476
rect 97692 140354 97748 140364
rect 96908 139048 96964 139244
rect 106652 139048 106708 155596
rect 106764 147140 106820 160076
rect 109340 148708 109396 160104
rect 112028 155540 112084 160104
rect 112028 155474 112084 155484
rect 109340 148642 109396 148652
rect 106764 147074 106820 147084
rect 112588 143780 112644 143790
rect 112588 142548 112644 143724
rect 114716 143780 114772 160104
rect 117404 157332 117460 160104
rect 117404 157266 117460 157276
rect 114716 143714 114772 143724
rect 116732 155764 116788 155774
rect 112588 139076 112644 142492
rect 114716 141204 114772 141214
rect 112588 139020 112952 139076
rect 114716 139048 114772 141148
rect 116732 139860 116788 155708
rect 118188 148708 118244 148718
rect 116732 139076 116788 139804
rect 116424 139020 116788 139076
rect 117516 147140 117572 147150
rect 117516 140868 117572 147084
rect 117516 139048 117572 140812
rect 118188 138740 118244 148652
rect 120092 147924 120148 160104
rect 120092 147858 120148 147868
rect 122668 160076 122808 160132
rect 122668 141428 122724 160076
rect 123564 157220 123620 157230
rect 119308 141204 119364 141214
rect 119308 139048 119364 141148
rect 122668 138852 122724 141372
rect 123340 147924 123396 147934
rect 123340 139076 123396 147868
rect 123564 141540 123620 157164
rect 123564 139076 123620 141484
rect 125020 145684 125076 145694
rect 124348 141316 124404 141326
rect 124348 140756 124404 141260
rect 124348 140690 124404 140700
rect 123564 139020 123816 139076
rect 125020 139048 125076 145628
rect 125468 140756 125524 160104
rect 128156 141988 128212 160104
rect 130872 160076 131012 160132
rect 128156 141922 128212 141932
rect 129276 142660 129332 142670
rect 129276 141988 129332 142604
rect 130956 142324 131012 160076
rect 133532 155652 133588 160104
rect 133532 155586 133588 155596
rect 133756 157332 133812 157342
rect 130956 142258 131012 142268
rect 133084 144116 133140 144126
rect 129276 141922 129332 141932
rect 125468 140690 125524 140700
rect 133084 139048 133140 144060
rect 133756 139636 133812 157276
rect 133756 139048 133812 139580
rect 133980 157108 134036 157118
rect 133980 141428 134036 157052
rect 133980 139076 134036 141372
rect 134652 155428 134708 155438
rect 134652 141876 134708 155372
rect 136220 145572 136276 160104
rect 138908 155764 138964 160104
rect 138908 155698 138964 155708
rect 141596 155428 141652 160104
rect 141596 155362 141652 155372
rect 144284 152068 144340 160104
rect 146972 159572 147028 160104
rect 146972 159506 147028 159516
rect 149100 157332 149156 157342
rect 144284 152002 144340 152012
rect 146972 157220 147028 157230
rect 136220 145506 136276 145516
rect 146972 145460 147028 157164
rect 146972 145394 147028 145404
rect 148428 148708 148484 148718
rect 143836 144452 143892 144462
rect 134652 139076 134708 141820
rect 133980 139020 134232 139076
rect 134568 139020 134708 139076
rect 134988 143780 135044 143790
rect 134988 139076 135044 143724
rect 135660 143780 135716 143790
rect 134988 139048 135492 139076
rect 135660 139048 135716 143724
rect 143836 139048 143892 144396
rect 144732 142772 144788 142782
rect 144732 139076 144788 142716
rect 135016 139020 135492 139048
rect 144648 139020 144788 139076
rect 145404 142436 145460 142446
rect 145404 141204 145460 142380
rect 145404 139048 145460 141148
rect 123340 139010 123396 139020
rect 122668 138786 122724 138796
rect 118188 138674 118244 138684
rect 135436 138628 135492 139020
rect 135436 138562 135492 138572
rect 142828 40292 142884 40302
rect 97020 39508 97076 39518
rect 72268 37940 72324 37950
rect 66556 4452 66612 4462
rect 60284 4162 60340 4172
rect 60844 4340 60900 4350
rect 60060 4050 60116 4060
rect 60844 480 60900 4284
rect 64652 4228 64708 4238
rect 62748 4116 62804 4126
rect 62748 480 62804 4060
rect 64652 480 64708 4172
rect 66556 480 66612 4396
rect 68684 4340 68740 4350
rect 68684 480 68740 4284
rect 49420 392 49672 480
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 480
rect 53228 392 53480 480
rect 53256 -960 53480 392
rect 55160 392 55412 480
rect 55160 -960 55384 392
rect 57064 -960 57288 480
rect 58940 392 59192 480
rect 60844 392 61096 480
rect 62748 392 63000 480
rect 64652 392 64904 480
rect 66556 392 66808 480
rect 58968 -960 59192 392
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 66584 -960 66808 392
rect 68488 392 68740 480
rect 70364 4228 70420 4238
rect 70364 480 70420 4172
rect 72268 480 72324 37884
rect 76076 37828 76132 37838
rect 74172 4116 74228 4126
rect 74172 480 74228 4060
rect 76076 480 76132 37772
rect 95116 36148 95172 36158
rect 83692 26068 83748 26078
rect 78204 4228 78260 4238
rect 78204 480 78260 4172
rect 80108 4228 80164 4238
rect 80108 480 80164 4172
rect 82012 4228 82068 4238
rect 82012 480 82068 4172
rect 70364 392 70616 480
rect 72268 392 72520 480
rect 74172 392 74424 480
rect 76076 392 76328 480
rect 68488 -960 68712 392
rect 70392 -960 70616 392
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 76104 -960 76328 392
rect 78008 392 78260 480
rect 79912 392 80164 480
rect 81816 392 82068 480
rect 83692 480 83748 26012
rect 87500 24388 87556 24398
rect 85820 4340 85876 4350
rect 85820 480 85876 4284
rect 83692 392 83944 480
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 83720 -960 83944 392
rect 85624 392 85876 480
rect 87500 480 87556 24332
rect 91308 15988 91364 15998
rect 89628 6020 89684 6030
rect 89628 480 89684 5964
rect 87500 392 87752 480
rect 85624 -960 85848 392
rect 87528 -960 87752 392
rect 89432 392 89684 480
rect 91308 480 91364 15932
rect 93436 7588 93492 7598
rect 93436 480 93492 7532
rect 91308 392 91560 480
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 392 93492 480
rect 95116 480 95172 36092
rect 97020 480 97076 39452
rect 106540 37940 106596 37950
rect 104636 12628 104692 12638
rect 99036 7700 99092 7710
rect 99036 480 99092 7644
rect 101052 5908 101108 5918
rect 101052 480 101108 5852
rect 102956 4228 103012 4238
rect 102956 480 103012 4172
rect 95116 392 95368 480
rect 97020 392 97272 480
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 480
rect 100856 392 101108 480
rect 102760 392 103012 480
rect 104636 480 104692 12572
rect 106540 480 106596 37884
rect 110348 37828 110404 37838
rect 108668 4228 108724 4238
rect 108668 480 108724 4172
rect 104636 392 104888 480
rect 106540 392 106792 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 392 108724 480
rect 110348 480 110404 37772
rect 119868 36260 119924 36270
rect 112476 4228 112532 4238
rect 112476 480 112532 4172
rect 114380 4228 114436 4238
rect 114380 480 114436 4172
rect 118188 4228 118244 4238
rect 116284 4116 116340 4126
rect 116284 480 116340 4060
rect 118188 480 118244 4172
rect 110348 392 110600 480
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 392 112532 480
rect 114184 392 114436 480
rect 116088 392 116340 480
rect 117992 392 118244 480
rect 119868 480 119924 36204
rect 139132 5124 139188 5134
rect 133420 4788 133476 4798
rect 121996 4676 122052 4686
rect 121996 480 122052 4620
rect 127596 4564 127652 4574
rect 125804 4452 125860 4462
rect 123900 4340 123956 4350
rect 123900 480 123956 4284
rect 125804 480 125860 4396
rect 127596 480 127652 4508
rect 131516 4116 131572 4126
rect 129612 4004 129668 4014
rect 129612 480 129668 3948
rect 131516 480 131572 4060
rect 133420 480 133476 4732
rect 135324 4676 135380 4686
rect 135324 480 135380 4620
rect 137228 3444 137284 3454
rect 137228 480 137284 3388
rect 139132 480 139188 5068
rect 141036 4900 141092 4910
rect 141036 480 141092 4844
rect 142828 480 142884 40236
rect 146748 5012 146804 5022
rect 144844 4788 144900 4798
rect 144844 480 144900 4732
rect 146748 480 146804 4956
rect 119868 392 120120 480
rect 112280 -960 112504 392
rect 114184 -960 114408 392
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 392 122052 480
rect 123704 392 123956 480
rect 125608 392 125860 480
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 480
rect 129416 392 129668 480
rect 131320 392 131572 480
rect 133224 392 133476 480
rect 135128 392 135380 480
rect 137032 392 137284 480
rect 138936 392 139188 480
rect 140840 392 141092 480
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144648 392 144900 480
rect 146552 392 146804 480
rect 148428 480 148484 148652
rect 148652 144004 148708 144014
rect 148652 4340 148708 143948
rect 148876 143892 148932 143902
rect 148876 4564 148932 143836
rect 149100 143668 149156 157276
rect 149660 144452 149716 160104
rect 149660 144386 149716 144396
rect 150332 147252 150388 147262
rect 149100 143602 149156 143612
rect 148876 4498 148932 4508
rect 148652 4274 148708 4284
rect 150332 480 150388 147196
rect 150444 145796 150500 145806
rect 150444 4452 150500 145740
rect 152012 145460 152068 145470
rect 152012 4788 152068 145404
rect 152348 143780 152404 160104
rect 153692 156324 153748 156334
rect 153692 144116 153748 156268
rect 155036 156324 155092 160104
rect 157276 158900 157332 158910
rect 155036 156258 155092 156268
rect 155372 157108 155428 157118
rect 153692 144050 153748 144060
rect 154140 144228 154196 144238
rect 152348 143714 152404 143724
rect 152572 143780 152628 143790
rect 152012 4722 152068 4732
rect 150444 4386 150500 4396
rect 152460 4340 152516 4350
rect 152460 480 152516 4284
rect 152572 4116 152628 143724
rect 152572 4050 152628 4060
rect 148428 392 148680 480
rect 150332 392 150584 480
rect 144648 -960 144872 392
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 392 152516 480
rect 154140 480 154196 144172
rect 155372 4676 155428 157052
rect 157276 4900 157332 158844
rect 157276 4834 157332 4844
rect 157500 147140 157556 147150
rect 155372 4610 155428 4620
rect 157500 4564 157556 147084
rect 157724 145684 157780 160104
rect 160412 157332 160468 160104
rect 160412 157266 160468 157276
rect 162092 156324 162148 156334
rect 160860 152404 160916 152414
rect 157724 145618 157780 145628
rect 159852 145684 159908 145694
rect 157500 4498 157556 4508
rect 157948 143668 158004 143678
rect 156156 4228 156212 4238
rect 156156 480 156212 4172
rect 157948 480 158004 143612
rect 159852 480 159908 145628
rect 160860 4676 160916 152348
rect 162092 147028 162148 156268
rect 163100 156324 163156 160104
rect 165788 157220 165844 160104
rect 165788 157154 165844 157164
rect 163100 156258 163156 156268
rect 168476 150388 168532 160104
rect 168476 150322 168532 150332
rect 162092 146962 162148 146972
rect 171164 147028 171220 160104
rect 173880 160076 174692 160132
rect 174636 156324 174692 160076
rect 174636 156268 174804 156324
rect 174748 150500 174804 156268
rect 174748 150434 174804 150444
rect 176092 152852 176148 152862
rect 171164 146962 171220 146972
rect 173516 145684 173572 145694
rect 165340 144116 165396 144126
rect 163772 142324 163828 142334
rect 163772 139048 163828 142268
rect 164556 142324 164612 142334
rect 164556 141988 164612 142268
rect 164556 141922 164612 141932
rect 164444 141316 164500 141326
rect 164444 139048 164500 141260
rect 165340 139048 165396 144060
rect 173516 139048 173572 145628
rect 174188 142660 174244 142670
rect 174188 139748 174244 142604
rect 174188 139048 174244 139692
rect 174636 142212 174692 142222
rect 174636 141652 174692 142156
rect 174636 139076 174692 141596
rect 174552 139020 174692 139076
rect 174972 142100 175028 142110
rect 174972 139048 175028 142044
rect 175420 140756 175476 140766
rect 175420 139076 175476 140700
rect 176092 139048 176148 152796
rect 176540 147140 176596 160104
rect 179228 157332 179284 160104
rect 179228 157266 179284 157276
rect 181916 147924 181972 160104
rect 184604 152852 184660 160104
rect 184604 152786 184660 152796
rect 181916 147858 181972 147868
rect 184268 147924 184324 147934
rect 176540 147074 176596 147084
rect 176316 142100 176372 142110
rect 176316 141764 176372 142044
rect 176316 141698 176372 141708
rect 184268 139048 184324 147868
rect 187292 145684 187348 160104
rect 187292 145618 187348 145628
rect 188972 156324 189028 156334
rect 188972 144116 189028 156268
rect 189980 156324 190036 160104
rect 192668 157108 192724 160104
rect 195356 157220 195412 160104
rect 198072 160076 198212 160132
rect 195356 157154 195412 157164
rect 192668 157042 192724 157052
rect 198156 156324 198212 160076
rect 198156 156268 198324 156324
rect 189980 156258 190036 156268
rect 198268 150612 198324 156268
rect 200732 155876 200788 160104
rect 200732 155810 200788 155820
rect 203420 152292 203476 160104
rect 203420 152226 203476 152236
rect 198268 150546 198324 150556
rect 188972 144050 189028 144060
rect 206108 144116 206164 160104
rect 208796 157444 208852 160104
rect 208796 157378 208852 157388
rect 211484 147364 211540 160104
rect 214172 155540 214228 160104
rect 216860 157556 216916 160104
rect 216860 157490 216916 157500
rect 214172 155474 214228 155484
rect 219548 150388 219604 160104
rect 222236 152180 222292 160104
rect 224952 160076 225092 160132
rect 222236 152114 222292 152124
rect 222572 157332 222628 157342
rect 219548 150322 219604 150332
rect 211484 147298 211540 147308
rect 206108 144050 206164 144060
rect 206556 145572 206612 145582
rect 186396 142100 186452 142110
rect 185052 141204 185108 141214
rect 185052 139048 185108 141148
rect 186396 141204 186452 142044
rect 186396 141138 186452 141148
rect 193340 140644 193396 140654
rect 192780 140532 192836 140542
rect 191996 140420 192052 140430
rect 190988 140308 191044 140318
rect 185724 140196 185780 140206
rect 185724 139076 185780 140140
rect 185612 139048 185780 139076
rect 190988 139972 191044 140252
rect 190988 139048 191044 139916
rect 191996 140084 192052 140364
rect 191996 139048 192052 140028
rect 192780 139524 192836 140476
rect 192780 139048 192836 139468
rect 193340 140308 193396 140588
rect 193340 139048 193396 140252
rect 196700 139188 196756 139198
rect 175420 139010 175476 139020
rect 185612 139020 185752 139048
rect 185612 138852 185668 139020
rect 196700 138852 196756 139132
rect 206556 139048 206612 145516
rect 222572 144004 222628 157276
rect 225036 156324 225092 160076
rect 225036 156268 225204 156324
rect 225148 153748 225204 156268
rect 225148 153682 225204 153692
rect 227612 145684 227668 160104
rect 230300 156548 230356 160104
rect 230300 156482 230356 156492
rect 232988 145796 233044 160104
rect 234332 156548 234388 156558
rect 232988 145730 233044 145740
rect 233100 147140 233156 147150
rect 227612 145618 227668 145628
rect 222572 143938 222628 143948
rect 224924 144004 224980 144014
rect 212940 142436 212996 142446
rect 212940 139048 212996 142380
rect 223804 141540 223860 141550
rect 214620 141204 214676 141214
rect 214620 139048 214676 141148
rect 219324 141204 219380 141214
rect 217420 140868 217476 140878
rect 216412 140532 216468 140542
rect 216412 139860 216468 140476
rect 216412 139048 216468 139804
rect 217420 140420 217476 140812
rect 217420 139048 217476 140364
rect 219324 139048 219380 141148
rect 223356 139412 223412 139422
rect 223356 138964 223412 139356
rect 223804 139048 223860 141484
rect 224924 139048 224980 143948
rect 233100 139048 233156 147084
rect 234332 144004 234388 156492
rect 234332 143938 234388 143948
rect 235676 143668 235732 160104
rect 235676 143602 235732 143612
rect 235788 150500 235844 150510
rect 235788 143444 235844 150444
rect 238364 145460 238420 160104
rect 241052 145572 241108 160104
rect 241948 157220 242004 157230
rect 241948 150724 242004 157164
rect 243740 156324 243796 160104
rect 246428 157220 246484 160104
rect 246428 157154 246484 157164
rect 247772 157444 247828 157454
rect 246652 157108 246708 157118
rect 243740 156258 243796 156268
rect 246092 156324 246148 156334
rect 241948 150658 242004 150668
rect 241052 145506 241108 145516
rect 243852 147028 243908 147038
rect 238364 145394 238420 145404
rect 235676 143388 235844 143444
rect 235004 142324 235060 142334
rect 234556 141876 234612 141886
rect 234220 141428 234276 141438
rect 233772 139636 233828 139646
rect 233772 139076 233828 139580
rect 233996 139188 234052 139198
rect 233996 139076 234052 139132
rect 233772 139048 234052 139076
rect 234220 139048 234276 141372
rect 234556 139048 234612 141820
rect 235004 141876 235060 142268
rect 235004 141810 235060 141820
rect 235116 142212 235172 142222
rect 235116 141428 235172 142156
rect 235116 141362 235172 141372
rect 235004 139300 235060 139310
rect 235004 139076 235060 139244
rect 234780 139048 235060 139076
rect 235676 139048 235732 143388
rect 243852 139048 243908 146972
rect 246092 143780 246148 156268
rect 246652 147252 246708 157052
rect 247772 147476 247828 157388
rect 249116 157108 249172 160104
rect 249116 157042 249172 157052
rect 251804 156324 251860 160104
rect 251804 156258 251860 156268
rect 252812 157556 252868 157566
rect 247772 147410 247828 147420
rect 249340 148708 249396 148718
rect 246652 147186 246708 147196
rect 246092 143714 246148 143724
rect 247548 146244 247604 146254
rect 244636 141204 244692 141214
rect 244636 139048 244692 141148
rect 245420 140644 245476 140654
rect 245420 139048 245476 140588
rect 233800 139020 234052 139048
rect 234780 139020 235032 139048
rect 223356 138898 223412 138908
rect 196924 138852 196980 138862
rect 196700 138796 196924 138852
rect 185612 138786 185668 138796
rect 196924 138786 196980 138796
rect 218204 138740 218260 138750
rect 218204 138674 218260 138684
rect 234780 138628 234836 139020
rect 234780 138562 234836 138572
rect 195916 39508 195972 39518
rect 176988 14308 177044 14318
rect 160860 4610 160916 4620
rect 175084 4676 175140 4686
rect 163884 4564 163940 4574
rect 161980 4452 162036 4462
rect 161980 480 162036 4396
rect 163884 480 163940 4508
rect 169596 4340 169652 4350
rect 167916 4228 167972 4238
rect 167692 4172 167916 4228
rect 165788 4116 165844 4126
rect 165788 480 165844 4060
rect 167692 480 167748 4172
rect 167916 4162 167972 4172
rect 169596 480 169652 4284
rect 171388 4228 171444 4238
rect 171388 480 171444 4172
rect 173404 3892 173460 3902
rect 173404 480 173460 3836
rect 154140 392 154392 480
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 480
rect 157948 392 158200 480
rect 159852 392 160104 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 392 162036 480
rect 163688 392 163940 480
rect 165592 392 165844 480
rect 167496 392 167748 480
rect 169400 392 169652 480
rect 161784 -960 162008 392
rect 163688 -960 163912 392
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 -960 171528 480
rect 173208 392 173460 480
rect 175084 480 175140 4620
rect 176988 480 177044 14252
rect 184604 12628 184660 12638
rect 182924 6132 182980 6142
rect 179116 4116 179172 4126
rect 179116 480 179172 4060
rect 181020 4116 181076 4126
rect 181020 480 181076 4060
rect 182924 480 182980 6076
rect 175084 392 175336 480
rect 176988 392 177240 480
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 392 179172 480
rect 180824 392 181076 480
rect 182728 392 182980 480
rect 184604 480 184660 12572
rect 186732 7700 186788 7710
rect 186732 480 186788 7644
rect 190540 7588 190596 7598
rect 188636 4116 188692 4126
rect 188636 480 188692 4060
rect 190540 480 190596 7532
rect 192444 4340 192500 4350
rect 192444 480 192500 4284
rect 194348 4228 194404 4238
rect 194348 480 194404 4172
rect 195916 4228 195972 39452
rect 197932 37940 197988 37950
rect 195916 4162 195972 4172
rect 196028 37828 196084 37838
rect 184604 392 184856 480
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 392
rect 186536 392 186788 480
rect 188440 392 188692 480
rect 190344 392 190596 480
rect 192248 392 192500 480
rect 194152 392 194404 480
rect 196028 480 196084 37772
rect 197932 480 197988 37884
rect 209356 36260 209412 36270
rect 201740 36148 201796 36158
rect 199948 29428 200004 29438
rect 199948 480 200004 29372
rect 201740 480 201796 36092
rect 207452 32788 207508 32798
rect 203644 31108 203700 31118
rect 203644 480 203700 31052
rect 205772 4452 205828 4462
rect 205772 480 205828 4396
rect 196028 392 196280 480
rect 197932 392 198184 480
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 392 205828 480
rect 207452 480 207508 32732
rect 209356 480 209412 36204
rect 221004 6020 221060 6030
rect 215292 5908 215348 5918
rect 211484 4564 211540 4574
rect 211484 480 211540 4508
rect 215292 480 215348 5852
rect 221004 480 221060 5964
rect 238140 4676 238196 4686
rect 226716 4116 226772 4126
rect 226716 480 226772 4060
rect 232428 4116 232484 4126
rect 232428 480 232484 4060
rect 238140 480 238196 4620
rect 247548 4340 247604 146188
rect 247548 4274 247604 4284
rect 243852 4228 243908 4238
rect 243852 480 243908 4172
rect 249340 480 249396 148652
rect 252812 147140 252868 157500
rect 254492 157332 254548 160104
rect 257180 159460 257236 160104
rect 259896 160076 260372 160132
rect 257180 159394 257236 159404
rect 260316 159012 260372 160076
rect 260316 158956 260484 159012
rect 260428 158900 260484 158956
rect 260428 158834 260484 158844
rect 262556 157892 262612 160104
rect 262556 157826 262612 157836
rect 265244 157556 265300 160104
rect 265244 157490 265300 157500
rect 254492 157266 254548 157276
rect 265468 157332 265524 157342
rect 261212 157220 261268 157230
rect 258636 156324 258692 156334
rect 258636 155652 258692 156268
rect 258636 155586 258692 155596
rect 252812 147074 252868 147084
rect 255052 152404 255108 152414
rect 250348 143892 250404 143902
rect 250348 4228 250404 143836
rect 250348 4162 250404 4172
rect 255052 480 255108 152348
rect 257852 151172 257908 151182
rect 257852 4564 257908 151116
rect 260316 148820 260372 148830
rect 257852 4498 257908 4508
rect 259532 138964 259588 138974
rect 259532 4452 259588 138908
rect 259532 4386 259588 4396
rect 260316 4228 260372 148764
rect 261212 143892 261268 157164
rect 264572 157108 264628 157118
rect 264572 147028 264628 157052
rect 265468 150500 265524 157276
rect 267932 157108 267988 160104
rect 270620 157780 270676 160104
rect 270620 157714 270676 157724
rect 273308 157668 273364 160104
rect 273868 158900 273924 158910
rect 273868 157892 273924 158844
rect 273868 157826 273924 157836
rect 275996 157892 276052 160104
rect 277676 159012 277732 300076
rect 277676 158946 277732 158956
rect 275996 157826 276052 157836
rect 273308 157602 273364 157612
rect 267932 157042 267988 157052
rect 265468 150434 265524 150444
rect 278796 148708 278852 305452
rect 278908 152404 278964 306796
rect 279020 160244 279076 309484
rect 279132 301476 279188 301486
rect 279132 160356 279188 301420
rect 284732 170548 284788 330988
rect 289772 266420 289828 373996
rect 294812 352548 294868 352558
rect 293132 324324 293188 324334
rect 289772 266354 289828 266364
rect 291452 322980 291508 322990
rect 284732 170482 284788 170492
rect 291452 162148 291508 322924
rect 293132 163828 293188 324268
rect 293132 163762 293188 163772
rect 291452 162082 291508 162092
rect 279132 160290 279188 160300
rect 279020 160178 279076 160188
rect 278908 152338 278964 152348
rect 278796 148642 278852 148652
rect 284284 152292 284340 152302
rect 273420 147476 273476 147486
rect 264572 146962 264628 146972
rect 265356 147364 265412 147374
rect 261212 143826 261268 143836
rect 263788 141988 263844 141998
rect 263788 138964 263844 141932
rect 264460 141876 264516 141886
rect 264460 141316 264516 141820
rect 264460 139048 264516 141260
rect 265356 139048 265412 147308
rect 273420 139048 273476 147420
rect 276108 144116 276164 144126
rect 274988 141764 275044 141774
rect 274540 141652 274596 141662
rect 274204 139748 274260 139758
rect 274204 139048 274260 139692
rect 274540 139048 274596 141596
rect 274988 141428 275044 141708
rect 274988 139048 275044 141372
rect 275436 139076 275492 139086
rect 263788 138898 263844 138908
rect 275324 139020 275436 139076
rect 276108 139048 276164 144060
rect 284284 139048 284340 152236
rect 294812 152292 294868 352492
rect 294924 264852 294980 375340
rect 296492 372708 296548 372718
rect 296492 273140 296548 372652
rect 388892 368788 388948 368798
rect 299852 353892 299908 353902
rect 296492 273074 296548 273084
rect 298172 329700 298228 329710
rect 294924 264786 294980 264796
rect 298172 168868 298228 329644
rect 299852 271684 299908 353836
rect 299852 271618 299908 271628
rect 303212 280028 303576 280084
rect 298172 168802 298228 168812
rect 294812 152226 294868 152236
rect 285068 142100 285124 142110
rect 285068 141316 285124 142044
rect 285068 139048 285124 141260
rect 303212 140644 303268 280028
rect 304220 275266 304276 280056
rect 304220 275214 304222 275266
rect 304274 275214 304276 275266
rect 304220 275202 304276 275214
rect 304444 280028 305032 280084
rect 304444 270004 304500 280028
rect 308252 275716 308308 275726
rect 304444 269938 304500 269948
rect 304892 275266 304948 275278
rect 304892 275214 304894 275266
rect 304946 275214 304948 275266
rect 304892 149548 304948 275214
rect 308252 216020 308308 275660
rect 308252 215954 308308 215964
rect 309932 275604 309988 275614
rect 309932 214340 309988 275548
rect 313292 275604 313348 280056
rect 313964 278908 314020 280056
rect 314328 280028 314580 280084
rect 314776 280028 315028 280084
rect 315224 280028 315700 280084
rect 314524 278908 314580 280028
rect 314972 278908 315028 280028
rect 315644 278908 315700 280028
rect 313964 278852 314132 278908
rect 314524 278852 314692 278908
rect 314972 278852 315588 278908
rect 315644 278852 315812 278908
rect 313292 275538 313348 275548
rect 309932 214274 309988 214284
rect 308252 157108 308308 157118
rect 308252 156212 308308 157052
rect 308252 156146 308308 156156
rect 304780 149492 304948 149548
rect 306572 155764 306628 155774
rect 304780 142772 304836 149492
rect 304780 142706 304836 142716
rect 303212 140578 303268 140588
rect 293356 140308 293412 140318
rect 285740 140196 285796 140206
rect 285740 139860 285796 140140
rect 292012 140084 292068 140094
rect 285740 139048 285796 139804
rect 291004 139972 291060 139982
rect 291004 139048 291060 139916
rect 292012 139636 292068 140028
rect 292012 139048 292068 139580
rect 292796 140084 292852 140094
rect 292796 139524 292852 140028
rect 292796 139048 292852 139468
rect 293356 139524 293412 140252
rect 293356 139048 293412 139468
rect 306572 139048 306628 155708
rect 312508 142996 312564 143006
rect 312508 139300 312564 142940
rect 314076 142996 314132 278852
rect 314636 273026 314692 278852
rect 314636 272974 314638 273026
rect 314690 272974 314692 273026
rect 314636 272962 314692 272974
rect 314076 142930 314132 142940
rect 315420 144116 315476 144126
rect 315420 143220 315476 144060
rect 312508 139234 312564 139244
rect 312956 142436 313012 142446
rect 312956 139048 313012 142380
rect 314636 141204 314692 141214
rect 314636 139048 314692 141148
rect 315420 139188 315476 143164
rect 315532 143332 315588 278852
rect 315532 142212 315588 143276
rect 315644 273026 315700 273038
rect 315644 272974 315646 273026
rect 315698 272974 315700 273026
rect 315644 143108 315700 272974
rect 315756 144116 315812 278852
rect 315868 275716 315924 280056
rect 315868 275650 315924 275660
rect 322588 280028 323960 280084
rect 322588 222740 322644 280028
rect 324380 273026 324436 273038
rect 324380 272974 324382 273026
rect 324434 272974 324436 273026
rect 324380 267148 324436 272974
rect 325164 267148 325220 280056
rect 325388 280028 325528 280084
rect 325388 273026 325444 280028
rect 329644 275604 329700 280056
rect 329644 275538 329700 275548
rect 325388 272974 325390 273026
rect 325442 272974 325444 273026
rect 325388 272962 325444 272974
rect 330764 267148 330820 280056
rect 331464 280028 332388 280084
rect 332332 278908 332388 280028
rect 332332 278852 332500 278908
rect 322588 222674 322644 222684
rect 324268 267092 324436 267148
rect 325052 267092 325220 267148
rect 330316 267092 330820 267148
rect 330876 276388 330932 276398
rect 330876 275604 330932 276332
rect 315756 144050 315812 144060
rect 315756 143108 315812 143118
rect 315644 143052 315756 143108
rect 315756 142324 315812 143052
rect 324268 142660 324324 267092
rect 323596 142604 324324 142660
rect 324940 155876 324996 155886
rect 315756 142258 315812 142268
rect 316428 142324 316484 142334
rect 315532 142146 315588 142156
rect 315420 139122 315476 139132
rect 316428 140532 316484 142268
rect 316428 139048 316484 140476
rect 317436 142100 317492 142110
rect 317436 140420 317492 142044
rect 317436 139048 317492 140364
rect 318220 141764 318276 141774
rect 318220 139076 318276 141708
rect 317772 139048 318276 139076
rect 319228 141204 319284 141214
rect 319228 139048 319284 141148
rect 323596 139300 323652 142604
rect 323596 139076 323652 139244
rect 275324 138628 275380 139020
rect 275436 139010 275492 139020
rect 317772 139020 318248 139048
rect 323400 139020 323652 139076
rect 323820 142436 323876 142446
rect 323820 141540 323876 142380
rect 323820 139048 323876 141484
rect 324940 139048 324996 155820
rect 325052 142436 325108 267092
rect 325052 142370 325108 142380
rect 330316 262724 330372 267092
rect 330316 141764 330372 262668
rect 330876 142772 330932 275548
rect 332444 262948 332500 278852
rect 330876 142706 330932 142716
rect 331772 262164 331828 262174
rect 331772 142324 331828 262108
rect 330316 141698 330372 141708
rect 330876 141764 330932 141774
rect 330876 139188 330932 141708
rect 331772 140980 331828 142268
rect 332444 142100 332500 262892
rect 332556 262164 332612 280056
rect 332556 262098 332612 262108
rect 333452 280028 334264 280084
rect 334572 280028 335944 280084
rect 342328 280028 342692 280084
rect 332444 142034 332500 142044
rect 333116 150612 333172 150622
rect 331772 140914 331828 140924
rect 330876 139122 330932 139132
rect 333116 139048 333172 150556
rect 333452 142772 333508 280028
rect 334572 267148 334628 280028
rect 334348 267092 334628 267148
rect 334124 143332 334180 143342
rect 333452 142706 333508 142716
rect 333788 143220 333844 143230
rect 296828 138852 296884 138862
rect 296828 138786 296884 138796
rect 317772 138740 317828 139020
rect 317772 138674 317828 138684
rect 333788 138740 333844 143164
rect 334124 141988 334180 143276
rect 334124 139048 334180 141932
rect 334348 142884 334404 267092
rect 342636 215908 342692 280028
rect 342636 215842 342692 215852
rect 347788 279860 347844 279870
rect 335692 150724 335748 150734
rect 334348 141764 334404 142828
rect 334348 141698 334404 141708
rect 334572 143108 334628 143118
rect 334572 141540 334628 143052
rect 334572 139048 334628 141484
rect 335020 142996 335076 143006
rect 335020 140644 335076 142940
rect 335020 139048 335076 140588
rect 335692 139048 335748 150668
rect 343868 147252 343924 147262
rect 336028 142100 336084 142110
rect 336028 140196 336084 142044
rect 336028 140130 336084 140140
rect 343868 139048 343924 147196
rect 344652 142100 344708 142110
rect 344652 139048 344708 142044
rect 345324 141204 345380 141214
rect 345324 139076 345380 141148
rect 345324 139010 345380 139020
rect 333788 138674 333844 138684
rect 275324 138562 275380 138572
rect 260316 4162 260372 4172
rect 260764 14308 260820 14318
rect 260764 480 260820 14252
rect 317884 7588 317940 7598
rect 295036 6020 295092 6030
rect 283612 5124 283668 5134
rect 266700 4340 266756 4350
rect 266700 480 266756 4284
rect 272188 4228 272244 4238
rect 272188 480 272244 4172
rect 277900 4228 277956 4238
rect 277900 480 277956 4172
rect 283612 480 283668 5068
rect 289324 5124 289380 5134
rect 289324 480 289380 5068
rect 295036 480 295092 5964
rect 312172 6020 312228 6030
rect 300748 5124 300804 5134
rect 300748 480 300804 5068
rect 306460 4228 306516 4238
rect 306460 480 306516 4172
rect 312172 480 312228 5964
rect 317884 480 317940 7532
rect 346668 4340 346724 4350
rect 323596 4228 323652 4238
rect 323596 480 323652 4172
rect 329308 4228 329364 4238
rect 329308 480 329364 4172
rect 335244 4228 335300 4238
rect 335244 480 335300 4172
rect 340956 4228 341012 4238
rect 340956 480 341012 4172
rect 346668 480 346724 4284
rect 347788 4228 347844 279804
rect 347900 278404 347956 278414
rect 347900 4564 347956 278348
rect 350252 276836 350308 276846
rect 347900 4498 347956 4508
rect 348012 273252 348068 273262
rect 348012 4340 348068 273196
rect 350252 212548 350308 276780
rect 350252 212482 350308 212492
rect 350476 276612 350532 276622
rect 350476 5012 350532 276556
rect 352044 275604 352100 280056
rect 355544 280028 356020 280084
rect 356216 280028 356804 280084
rect 357000 280028 357812 280084
rect 358008 280028 359492 280084
rect 355292 279748 355348 279758
rect 352044 275538 352100 275548
rect 353948 275604 354004 275614
rect 353612 269892 353668 269902
rect 350476 4946 350532 4956
rect 352156 168868 352212 168878
rect 348012 4274 348068 4284
rect 347788 4162 347844 4172
rect 352156 480 352212 168812
rect 353612 20356 353668 269836
rect 353948 269892 354004 275548
rect 353948 269826 354004 269836
rect 353612 20290 353668 20300
rect 355292 4900 355348 279692
rect 355964 278908 356020 280028
rect 355964 278852 356132 278908
rect 356076 266644 356132 278852
rect 356748 268324 356804 280028
rect 356748 268258 356804 268268
rect 356076 266578 356132 266588
rect 357756 265076 357812 280028
rect 359436 270004 359492 280028
rect 363132 273252 363188 280056
rect 363804 275604 363860 280056
rect 363804 275538 363860 275548
rect 363132 273186 363188 273196
rect 359436 269938 359492 269948
rect 364588 268212 364644 280056
rect 371308 280028 372904 280084
rect 373464 280028 373716 280084
rect 373912 280028 374164 280084
rect 364588 268146 364644 268156
rect 366268 275604 366324 275614
rect 366268 268212 366324 275548
rect 366268 268146 366324 268156
rect 364476 266756 364532 266766
rect 357756 265010 357812 265020
rect 363804 265188 363860 265198
rect 357084 262836 357140 262846
rect 355292 4834 355348 4844
rect 356972 257908 357028 257918
rect 356972 4116 357028 257852
rect 357084 217700 357140 262780
rect 360332 262500 360388 262510
rect 360332 254548 360388 262444
rect 363804 259140 363860 265132
rect 364252 259140 364308 259150
rect 363804 259112 364252 259140
rect 363832 259084 364252 259112
rect 364252 259074 364308 259084
rect 364476 258804 364532 266700
rect 371308 266532 371364 280028
rect 373660 273026 373716 280028
rect 374108 278852 374164 280028
rect 374108 278786 374164 278796
rect 374332 273140 374388 280056
rect 374668 280028 374808 280084
rect 373660 272974 373662 273026
rect 373714 272974 373716 273026
rect 373660 272962 373716 272974
rect 373772 273084 374388 273140
rect 374444 278852 374500 278862
rect 371308 266466 371364 266476
rect 365372 262836 365428 262846
rect 365372 259112 365428 262780
rect 373772 262836 373828 273084
rect 374444 267148 374500 278796
rect 373772 262770 373828 262780
rect 374332 267092 374500 267148
rect 374556 273026 374612 273038
rect 374556 272974 374558 273026
rect 374610 272974 374612 273026
rect 373436 262500 373492 262510
rect 373436 259112 373492 262444
rect 374332 262500 374388 267092
rect 374556 263060 374612 272974
rect 374556 262994 374612 263004
rect 374332 262434 374388 262444
rect 374556 262836 374612 262846
rect 374220 262276 374276 262286
rect 374220 259140 374276 262220
rect 373884 259112 374276 259140
rect 373884 259084 374248 259112
rect 373884 259028 373940 259084
rect 373884 258962 373940 258972
rect 374556 258804 374612 262780
rect 374668 262276 374724 280028
rect 375452 276836 375508 280056
rect 375452 276770 375508 276780
rect 380492 275716 380548 275726
rect 380492 266756 380548 275660
rect 380492 266690 380548 266700
rect 382172 275604 382228 275614
rect 382172 264964 382228 275548
rect 383516 275604 383572 280056
rect 384412 275716 384468 280056
rect 384412 275650 384468 275660
rect 383516 275538 383572 275548
rect 383852 275604 383908 275614
rect 383852 265188 383908 275548
rect 385196 275604 385252 280056
rect 385196 275538 385252 275548
rect 385308 273252 385364 273262
rect 383852 265122 383908 265132
rect 385084 268212 385140 268222
rect 382172 264898 382228 264908
rect 375452 263060 375508 263070
rect 374668 262210 374724 262220
rect 375004 262500 375060 262510
rect 375004 259140 375060 262444
rect 375452 259140 375508 263004
rect 375004 259074 375060 259084
rect 375228 259112 375508 259140
rect 376124 262164 376180 262174
rect 376124 259112 376180 262108
rect 375228 259084 375480 259112
rect 363916 258776 364532 258804
rect 374332 258776 374612 258804
rect 363916 258748 364504 258776
rect 374332 258748 374584 258776
rect 363916 258692 363972 258748
rect 363916 258626 363972 258636
rect 374332 258692 374388 258748
rect 374332 258626 374388 258636
rect 375228 258692 375284 259084
rect 384300 258916 384356 258926
rect 385084 258916 385140 268156
rect 385308 259140 385364 273196
rect 388892 262612 388948 368732
rect 419132 342804 419188 342814
rect 419132 302428 419188 342748
rect 419132 302372 419412 302428
rect 419356 276388 419412 302372
rect 456092 276724 456148 429996
rect 460236 418180 460292 418190
rect 460124 416612 460180 416622
rect 456092 276658 456148 276668
rect 459452 381444 459508 381454
rect 388892 262546 388948 262556
rect 390572 270004 390628 270014
rect 385756 259140 385812 259150
rect 385308 259084 385756 259140
rect 385756 259074 385812 259084
rect 390572 259140 390628 269948
rect 396844 269892 396900 269902
rect 392812 268324 392868 268334
rect 391916 265076 391972 265086
rect 391916 259140 391972 265020
rect 392812 259140 392868 268268
rect 390628 259084 391048 259140
rect 391916 259112 392308 259140
rect 391944 259084 392308 259112
rect 390572 259046 390628 259084
rect 392252 259028 392308 259084
rect 392252 258962 392308 258972
rect 392476 259112 392868 259140
rect 393372 266644 393428 266654
rect 393372 259140 393428 266588
rect 393932 259140 393988 259150
rect 393372 259112 393932 259140
rect 392476 259084 392840 259112
rect 393400 259084 393932 259112
rect 396844 259140 396900 269836
rect 417452 262948 417508 262958
rect 416332 262388 416388 262398
rect 397292 259140 397348 259150
rect 396844 259112 397292 259140
rect 396872 259084 397292 259112
rect 416332 259112 416388 262332
rect 417452 259112 417508 262892
rect 418124 262724 418180 262734
rect 418124 259112 418180 262668
rect 419356 259140 419412 276332
rect 454972 271684 455028 271694
rect 423948 261380 424004 261390
rect 424004 261324 424228 261380
rect 423948 261314 424004 261324
rect 419272 259084 419412 259140
rect 424172 259140 424228 261324
rect 435708 260484 435764 260494
rect 432236 259812 432292 259822
rect 432236 259140 432292 259756
rect 424172 259084 424984 259140
rect 432236 259084 433048 259140
rect 435708 259112 435764 260428
rect 443436 259700 443492 259710
rect 443436 259140 443492 259644
rect 443436 259084 443912 259140
rect 392476 259028 392532 259084
rect 393932 259074 393988 259084
rect 397292 259074 397348 259084
rect 392476 258962 392532 258972
rect 385420 258916 385476 258926
rect 385084 258888 385420 258916
rect 385112 258860 385420 258888
rect 384300 258850 384356 258860
rect 385420 258850 385476 258860
rect 406588 258804 406644 258814
rect 406588 258738 406644 258748
rect 412412 258804 412468 258814
rect 414092 258804 414148 258814
rect 424396 258804 424452 258814
rect 412468 258748 413000 258804
rect 414148 258748 414680 258804
rect 423752 258748 424396 258804
rect 412412 258738 412468 258748
rect 414092 258738 414148 258748
rect 424396 258738 424452 258748
rect 375228 258626 375284 258636
rect 434924 258692 434980 258702
rect 434924 258626 434980 258636
rect 433804 258580 433860 258590
rect 433804 258514 433860 258524
rect 423388 258468 423444 258478
rect 423388 258402 423444 258412
rect 434140 258468 434196 258478
rect 434140 258402 434196 258412
rect 434588 258468 434644 258478
rect 434588 258402 434644 258412
rect 444668 258468 444724 258478
rect 444668 258402 444724 258412
rect 445340 258468 445396 258478
rect 445340 258402 445396 258412
rect 360332 254482 360388 254492
rect 357084 217634 357140 217644
rect 356972 4050 357028 4060
rect 357868 170548 357924 170558
rect 357868 480 357924 170492
rect 443884 155540 443940 155550
rect 406588 155428 406644 155438
rect 384412 153748 384468 153758
rect 365372 145796 365428 145806
rect 364252 142324 364308 142334
rect 364252 139076 364308 142268
rect 363832 139048 364308 139076
rect 364476 142324 364532 142334
rect 364476 141876 364532 142268
rect 364476 139048 364532 141820
rect 365372 139048 365428 145740
rect 376124 145684 376180 145694
rect 373436 144004 373492 144014
rect 373324 141876 373380 141886
rect 373324 141428 373380 141820
rect 373324 141362 373380 141372
rect 373436 139048 373492 143948
rect 374556 142212 374612 142222
rect 374556 141204 374612 142156
rect 374220 139748 374276 139758
rect 374220 139048 374276 139692
rect 374556 139048 374612 141148
rect 375004 141876 375060 141886
rect 375004 139048 375060 141820
rect 375452 141428 375508 141438
rect 375452 139076 375508 141372
rect 375228 139048 375508 139076
rect 376124 139048 376180 145628
rect 384412 139076 384468 153692
rect 363804 139020 364308 139048
rect 375228 139020 375480 139048
rect 384328 139020 384468 139076
rect 385084 141316 385140 141326
rect 385084 139048 385140 141260
rect 391916 140868 391972 140878
rect 391020 140308 391076 140318
rect 391020 139972 391076 140252
rect 385756 139860 385812 139870
rect 385756 139048 385812 139804
rect 391020 139048 391076 139916
rect 391916 139636 391972 140812
rect 393372 140756 393428 140766
rect 391916 139048 391972 139580
rect 392812 140532 392868 140542
rect 392812 140084 392868 140476
rect 392812 139048 392868 140028
rect 393372 139524 393428 140700
rect 393372 139048 393428 139468
rect 406588 139048 406644 155372
rect 424956 152180 425012 152190
rect 412412 142772 412468 142782
rect 412412 141764 412468 142716
rect 412412 139076 412468 141708
rect 423724 142436 423780 142446
rect 423724 141876 423780 142380
rect 414652 141204 414708 141214
rect 412412 139020 413000 139076
rect 414652 139048 414708 141148
rect 419244 141204 419300 141214
rect 416332 140980 416388 140990
rect 416332 139048 416388 140924
rect 417452 140196 417508 140206
rect 417452 139048 417508 140140
rect 417676 139188 417732 139198
rect 417676 139076 417732 139132
rect 417676 139048 418152 139076
rect 419244 139048 419300 141148
rect 423612 139188 423668 139198
rect 423612 139076 423668 139132
rect 417676 139020 418180 139048
rect 423416 139020 423668 139076
rect 423724 139048 423780 141820
rect 424956 139048 425012 152124
rect 433132 150388 433188 150398
rect 433132 139076 433188 150332
rect 435708 147140 435764 147150
rect 434140 141988 434196 141998
rect 433048 139020 433188 139076
rect 433804 141764 433860 141774
rect 433804 140084 433860 141708
rect 363804 138964 363860 139020
rect 363804 138898 363860 138908
rect 375228 138628 375284 139020
rect 418124 138964 418180 139020
rect 418124 138898 418180 138908
rect 396844 138852 396900 138862
rect 396844 138786 396900 138796
rect 433804 138740 433860 140028
rect 434140 139048 434196 141932
rect 434588 141540 434644 141550
rect 434588 139048 434644 141484
rect 434812 140644 434868 140654
rect 434812 138740 434868 140588
rect 435708 139048 435764 147084
rect 443884 139048 443940 155484
rect 449260 152292 449316 152302
rect 444668 141988 444724 141998
rect 444668 139048 444724 141932
rect 445564 139076 445620 139086
rect 445368 139020 445564 139076
rect 445564 139010 445620 139020
rect 434924 138740 434980 138750
rect 434812 138684 434924 138740
rect 433804 138674 433860 138684
rect 434924 138674 434980 138684
rect 375228 138562 375284 138572
rect 437836 36148 437892 36158
rect 426412 17668 426468 17678
rect 420700 15988 420756 15998
rect 392140 14308 392196 14318
rect 363580 5012 363636 5022
rect 363580 480 363636 4956
rect 375004 4900 375060 4910
rect 369292 4116 369348 4126
rect 369292 480 369348 4060
rect 375004 480 375060 4844
rect 380716 4788 380772 4798
rect 380716 480 380772 4732
rect 386428 4676 386484 4686
rect 386428 480 386484 4620
rect 392140 480 392196 14252
rect 409276 5908 409332 5918
rect 403564 4564 403620 4574
rect 397852 4452 397908 4462
rect 397852 480 397908 4396
rect 403564 480 403620 4508
rect 409276 480 409332 5852
rect 414988 4340 415044 4350
rect 414988 480 415044 4284
rect 420700 480 420756 15932
rect 426412 480 426468 17612
rect 432124 4228 432180 4238
rect 432124 480 432180 4172
rect 437836 480 437892 36092
rect 443772 4228 443828 4238
rect 443772 480 443828 4172
rect 449260 480 449316 152236
rect 454972 480 455028 271628
rect 459452 4228 459508 381388
rect 460124 37828 460180 416556
rect 460124 37762 460180 37772
rect 460236 36148 460292 418124
rect 461132 377860 461188 565292
rect 461244 432740 461300 570332
rect 462812 432852 462868 588924
rect 462812 432786 462868 432796
rect 462924 555268 462980 555278
rect 461244 432674 461300 432684
rect 461132 377794 461188 377804
rect 462812 430164 462868 430174
rect 462812 149716 462868 430108
rect 462924 377748 462980 555212
rect 464492 444500 464548 591276
rect 474348 583828 474404 595560
rect 474348 583762 474404 583772
rect 496412 582260 496468 595560
rect 518476 590996 518532 595560
rect 518476 590930 518532 590940
rect 496412 582194 496468 582204
rect 540540 582148 540596 595560
rect 540540 582082 540596 582092
rect 562604 578788 562660 595560
rect 584668 591332 584724 595560
rect 584668 591266 584724 591276
rect 562604 578722 562660 578732
rect 464492 444434 464548 444444
rect 464604 555380 464660 555390
rect 464604 432964 464660 555324
rect 468524 551572 468580 551582
rect 468412 551460 468468 551470
rect 468300 551348 468356 551358
rect 468188 551236 468244 551246
rect 467740 549556 467796 549566
rect 467740 501620 467796 549500
rect 468076 549108 468132 549118
rect 467740 501554 467796 501564
rect 467852 548324 467908 548334
rect 467740 495572 467796 495582
rect 467740 450436 467796 495516
rect 467852 453236 467908 548268
rect 467964 546980 468020 546990
rect 467964 459284 468020 546924
rect 468076 465332 468132 549052
rect 468076 465266 468132 465276
rect 468188 507668 468244 551180
rect 467964 459218 468020 459228
rect 467852 453170 467908 453180
rect 467740 450370 467796 450380
rect 464604 432898 464660 432908
rect 468188 393092 468244 507612
rect 468300 513716 468356 551292
rect 468300 394660 468356 513660
rect 468412 519764 468468 551404
rect 468412 396228 468468 519708
rect 468524 525812 468580 551516
rect 468524 397796 468580 525756
rect 468636 549444 468692 549454
rect 468636 531860 468692 549388
rect 495516 537796 495572 537806
rect 468636 446852 468692 531804
rect 470316 537684 470372 537694
rect 470092 500948 470148 500958
rect 468636 446786 468692 446796
rect 469868 459284 469924 459294
rect 468524 397730 468580 397740
rect 468636 421316 468692 421326
rect 468412 396162 468468 396172
rect 468300 394594 468356 394604
rect 468188 393026 468244 393036
rect 462924 377682 462980 377692
rect 467852 377188 467908 377198
rect 467852 160692 467908 377132
rect 467852 160626 467908 160636
rect 468636 159012 468692 421260
rect 469868 383684 469924 459228
rect 469980 403396 470036 403406
rect 469980 386820 470036 403340
rect 470092 391524 470148 500892
rect 470092 391458 470148 391468
rect 470204 464660 470260 464670
rect 469980 386754 470036 386764
rect 470204 385252 470260 464604
rect 470316 451556 470372 537628
rect 477596 537684 477652 537694
rect 477596 537572 477764 537628
rect 477708 534996 477764 537572
rect 495516 534996 495572 537740
rect 547148 537684 547204 537694
rect 512316 536004 512372 536014
rect 477708 534940 478296 534996
rect 495320 534940 495572 534996
rect 512204 535948 512316 536004
rect 512204 534996 512260 535948
rect 512316 535938 512372 535948
rect 547148 534996 547204 537628
rect 512204 534940 512344 534996
rect 546392 534940 547204 534996
rect 554428 537684 554484 537694
rect 529340 534324 529396 534334
rect 529340 534258 529396 534268
rect 470316 451490 470372 451500
rect 470652 452452 470708 452462
rect 470204 385186 470260 385196
rect 469868 383618 469924 383628
rect 470652 382116 470708 452396
rect 474908 450548 474964 450558
rect 474712 450492 474908 450548
rect 470876 450436 470932 450446
rect 470876 389956 470932 450380
rect 470876 389890 470932 389900
rect 472892 450324 472948 450334
rect 472892 388388 472948 450268
rect 474908 448420 474964 450492
rect 533036 450212 533092 450222
rect 474908 448354 474964 448364
rect 479612 448420 479668 448430
rect 477932 447972 477988 447982
rect 475132 447748 475188 447758
rect 474572 446852 474628 446862
rect 474572 399364 474628 446796
rect 474572 399298 474628 399308
rect 475132 398132 475188 447692
rect 477596 429828 477652 429838
rect 477036 422884 477092 422894
rect 476924 419748 476980 419758
rect 476252 415044 476308 415054
rect 476252 402948 476308 414988
rect 476252 402882 476308 402892
rect 476476 413476 476532 413486
rect 476476 402836 476532 413420
rect 476476 402770 476532 402780
rect 475132 398066 475188 398076
rect 472892 388322 472948 388332
rect 476252 397348 476308 397358
rect 470652 382050 470708 382060
rect 476252 334852 476308 397292
rect 476252 334786 476308 334796
rect 476364 383908 476420 383918
rect 476364 333956 476420 383852
rect 476924 379092 476980 419692
rect 476924 379026 476980 379036
rect 477036 375508 477092 422828
rect 477596 402276 477652 429772
rect 477596 402210 477652 402220
rect 477820 429716 477876 429726
rect 477820 399700 477876 429660
rect 477932 401492 477988 447916
rect 478492 447860 478548 447870
rect 478044 443268 478100 443278
rect 478044 402388 478100 443212
rect 478380 432068 478436 432078
rect 478044 402322 478100 402332
rect 478156 431956 478212 431966
rect 477932 401426 477988 401436
rect 478156 401380 478212 431900
rect 478380 402612 478436 432012
rect 478380 402546 478436 402556
rect 478156 401314 478212 401324
rect 478492 399812 478548 447804
rect 478716 426020 478772 426030
rect 478492 399746 478548 399756
rect 478604 424452 478660 424462
rect 477820 399634 477876 399644
rect 477036 375442 477092 375452
rect 477932 377412 477988 377422
rect 476364 333890 476420 333900
rect 476476 325892 476532 325902
rect 476252 324996 476308 325006
rect 476140 312452 476196 312462
rect 476140 293972 476196 312396
rect 476140 293906 476196 293916
rect 476252 292292 476308 324940
rect 476364 322308 476420 322318
rect 476364 297220 476420 322252
rect 476476 300580 476532 325836
rect 476700 324100 476756 324110
rect 476476 300514 476532 300524
rect 476588 314244 476644 314254
rect 476364 297154 476420 297164
rect 476252 292226 476308 292236
rect 476588 290612 476644 314188
rect 476700 300692 476756 324044
rect 476924 323204 476980 323214
rect 476700 300626 476756 300636
rect 476812 316932 476868 316942
rect 476812 297332 476868 316876
rect 476924 302372 476980 323148
rect 476924 302306 476980 302316
rect 477036 316036 477092 316046
rect 476812 297266 476868 297276
rect 476588 290546 476644 290556
rect 477036 289044 477092 315980
rect 477036 288978 477092 288988
rect 477932 266308 477988 377356
rect 478604 373828 478660 424396
rect 478604 373762 478660 373772
rect 478716 372148 478772 425964
rect 479612 379428 479668 448364
rect 480620 446964 480676 446974
rect 479612 379362 479668 379372
rect 480060 426916 480116 426926
rect 478716 372082 478772 372092
rect 479612 377300 479668 377310
rect 479612 271572 479668 377244
rect 480060 368900 480116 426860
rect 480620 400260 480676 446908
rect 484092 446964 484148 450072
rect 484092 446898 484148 446908
rect 488124 449652 488180 449662
rect 482748 444500 482804 444510
rect 482748 429912 482804 444444
rect 485436 432964 485492 432974
rect 484092 432852 484148 432862
rect 484092 429912 484148 432796
rect 485436 429912 485492 432908
rect 486780 432740 486836 432750
rect 486780 429912 486836 432684
rect 488124 429912 488180 449596
rect 493500 447972 493556 450072
rect 493500 447906 493556 447916
rect 502908 447860 502964 450072
rect 502908 447794 502964 447804
rect 504252 449540 504308 449550
rect 489468 437892 489524 437902
rect 489468 429912 489524 437836
rect 490812 432628 490868 432638
rect 490812 429912 490868 432572
rect 497532 432292 497588 432302
rect 496188 432180 496244 432190
rect 492156 432068 492212 432078
rect 492156 429912 492212 432012
rect 494844 431956 494900 431966
rect 493500 431844 493556 431854
rect 493500 429912 493556 431788
rect 494844 429912 494900 431900
rect 496188 429912 496244 432124
rect 497532 429912 497588 432236
rect 498876 432180 498932 432190
rect 498876 429912 498932 432124
rect 502908 432068 502964 432078
rect 502908 429912 502964 432012
rect 504252 429912 504308 449484
rect 512316 447748 512372 450072
rect 512316 447682 512372 447692
rect 521612 450044 521752 450100
rect 521612 448532 521668 450044
rect 521612 447412 521668 448476
rect 527436 449428 527492 449438
rect 527436 448532 527492 449372
rect 527436 448466 527492 448476
rect 531132 448532 531188 450072
rect 531132 448466 531188 448476
rect 521612 447346 521668 447356
rect 525756 447860 525812 447870
rect 509628 446180 509684 446190
rect 506940 444388 506996 444398
rect 505596 434420 505652 434430
rect 505596 429912 505652 434364
rect 506940 429912 506996 444332
rect 508284 437780 508340 437790
rect 508284 429912 508340 437724
rect 509628 429912 509684 446124
rect 510972 434308 511028 434318
rect 510972 429912 511028 434252
rect 512316 432628 512372 432638
rect 512316 429912 512372 432572
rect 519036 431956 519092 431966
rect 513660 429940 513716 429950
rect 519036 429912 519092 431900
rect 523068 431844 523124 431854
rect 521724 430276 521780 430286
rect 519596 430052 519652 430062
rect 519596 429940 519652 429996
rect 519596 429884 520408 429940
rect 521724 429912 521780 430220
rect 523068 429912 523124 431788
rect 524412 430164 524468 430174
rect 524412 429912 524468 430108
rect 525756 429912 525812 447804
rect 527100 447748 527156 447758
rect 527100 429912 527156 447692
rect 532700 446068 532756 446078
rect 532588 439348 532644 439358
rect 513660 429874 513716 429884
rect 515004 429828 515060 429838
rect 515004 429762 515060 429772
rect 516348 429716 516404 429726
rect 516348 429650 516404 429660
rect 517692 429492 517748 429502
rect 517692 429426 517748 429436
rect 500220 429380 500276 429390
rect 500220 429314 500276 429324
rect 501564 429268 501620 429278
rect 501564 429202 501620 429212
rect 532588 426468 532644 439292
rect 532588 426402 532644 426412
rect 532700 421092 532756 446012
rect 532700 421026 532756 421036
rect 532812 437668 532868 437678
rect 532812 415716 532868 437612
rect 532812 415650 532868 415660
rect 532924 429604 532980 429614
rect 532924 410340 532980 429548
rect 532924 410274 532980 410284
rect 480620 400194 480676 400204
rect 533036 383460 533092 450156
rect 540540 447860 540596 450072
rect 540540 447794 540596 447804
rect 549948 447748 550004 450072
rect 549948 447682 550004 447692
rect 533372 407428 533428 407438
rect 533372 404964 533428 407372
rect 554428 407428 554484 537628
rect 557788 508340 557844 508350
rect 557788 451332 557844 508284
rect 557788 451266 557844 451276
rect 557900 497812 557956 497822
rect 557900 451220 557956 497756
rect 557900 451154 557956 451164
rect 558012 487284 558068 487294
rect 558012 450324 558068 487228
rect 590492 482916 590548 482926
rect 558124 476756 558180 476766
rect 558124 451444 558180 476700
rect 558124 451378 558180 451388
rect 558236 466228 558292 466238
rect 558236 451108 558292 466172
rect 558236 451042 558292 451052
rect 590492 450548 590548 482860
rect 590492 450482 590548 450492
rect 558012 450258 558068 450268
rect 554428 407362 554484 407372
rect 533372 404898 533428 404908
rect 533372 390628 533428 390638
rect 533372 388836 533428 390572
rect 533372 388770 533428 388780
rect 533036 383394 533092 383404
rect 484764 380772 484820 380782
rect 484764 380706 484820 380716
rect 590604 380548 590660 380558
rect 502908 380436 502964 380446
rect 502908 380370 502964 380380
rect 526316 380436 526372 380446
rect 526372 380380 527128 380436
rect 526316 380370 526372 380380
rect 500892 380324 500948 380334
rect 500892 380258 500948 380268
rect 482748 380212 482804 380222
rect 482748 380146 482804 380156
rect 492828 380100 492884 380110
rect 486780 377748 486836 380072
rect 488796 377860 488852 380072
rect 488796 377794 488852 377804
rect 486780 377682 486836 377692
rect 490812 377636 490868 380072
rect 523068 380100 523124 380110
rect 492828 380034 492884 380044
rect 494844 377972 494900 380072
rect 496860 379540 496916 380072
rect 496860 379474 496916 379484
rect 494844 377906 494900 377916
rect 498876 377972 498932 380072
rect 498876 377906 498932 377916
rect 490812 377570 490868 377580
rect 504924 377524 504980 380072
rect 504924 377458 504980 377468
rect 480060 368834 480116 368844
rect 506940 368788 506996 380072
rect 508956 377412 509012 380072
rect 508956 377346 509012 377356
rect 510972 377300 511028 380072
rect 510972 377234 511028 377244
rect 512988 377188 513044 380072
rect 515004 379428 515060 380072
rect 515004 379362 515060 379372
rect 517020 378980 517076 380072
rect 519036 379652 519092 380072
rect 519036 379586 519092 379596
rect 517020 378914 517076 378924
rect 521052 377972 521108 380072
rect 523068 380034 523124 380044
rect 521052 377906 521108 377916
rect 525084 377972 525140 380072
rect 525084 377906 525140 377916
rect 559468 379092 559524 379102
rect 512988 377122 513044 377132
rect 506940 368722 506996 368732
rect 482524 348628 482580 348638
rect 482524 342804 482580 348572
rect 498988 345380 499044 345390
rect 495964 344932 496020 344942
rect 492604 344708 492660 344718
rect 482524 341880 482580 342748
rect 485884 344596 485940 344606
rect 485884 341880 485940 344540
rect 489244 344484 489300 344494
rect 489244 341880 489300 344428
rect 492604 341880 492660 344652
rect 495964 341880 496020 344876
rect 498988 341908 499044 345324
rect 502348 345380 502404 345390
rect 502348 341908 502404 345324
rect 505708 345380 505764 345390
rect 505708 341908 505764 345324
rect 509404 344484 509460 344494
rect 498988 341852 499352 341908
rect 502348 341852 502712 341908
rect 505708 341852 506072 341908
rect 509404 341880 509460 344428
rect 512764 344484 512820 344494
rect 512764 341880 512820 344428
rect 516124 344484 516180 344494
rect 516124 341880 516180 344428
rect 519484 344484 519540 344494
rect 519484 341880 519540 344428
rect 479612 271506 479668 271516
rect 477932 266242 477988 266252
rect 501228 160132 501284 160142
rect 468636 158946 468692 158956
rect 472892 160076 473592 160132
rect 474264 160076 474628 160132
rect 464716 155428 464772 155438
rect 462812 149650 462868 149660
rect 464492 150388 464548 150398
rect 463820 142772 463876 142782
rect 463820 142100 463876 142716
rect 463820 139048 463876 142044
rect 464492 142324 464548 150332
rect 464716 142772 464772 155372
rect 464716 142706 464772 142716
rect 465388 150500 465444 150510
rect 464492 139048 464548 142268
rect 465388 139048 465444 150444
rect 472892 141988 472948 160076
rect 474572 156324 474628 160076
rect 475020 159460 475076 160104
rect 475020 159394 475076 159404
rect 483196 158788 483252 160104
rect 483980 159684 484036 160104
rect 483980 159618 484036 159628
rect 484092 160076 484344 160132
rect 483196 158722 483252 158732
rect 474572 156258 474628 156268
rect 472892 141922 472948 141932
rect 473452 155652 473508 155662
rect 473452 139048 473508 155596
rect 474572 152180 474628 152190
rect 474124 147140 474180 147150
rect 474124 141204 474180 147084
rect 474124 139048 474180 141148
rect 474572 142212 474628 152124
rect 475468 150500 475524 150510
rect 474572 139048 474628 142156
rect 475020 145684 475076 145694
rect 475020 142548 475076 145628
rect 475020 139048 475076 142492
rect 475468 138740 475524 150444
rect 476028 147028 476084 147038
rect 476028 139048 476084 146972
rect 484092 141764 484148 160076
rect 484764 154868 484820 160104
rect 484652 154812 484820 154868
rect 484988 160076 485128 160132
rect 484092 141698 484148 141708
rect 484316 143892 484372 143902
rect 484316 139048 484372 143836
rect 484652 142100 484708 154812
rect 484988 149548 485044 160076
rect 485212 159684 485268 159694
rect 485268 159628 485492 159684
rect 485212 159618 485268 159628
rect 484652 142034 484708 142044
rect 484764 149492 485044 149548
rect 484764 140644 484820 149492
rect 485100 143892 485156 143902
rect 485100 142660 485156 143836
rect 484764 140084 484820 140588
rect 484764 140018 484820 140028
rect 484876 141764 484932 141774
rect 475244 138712 475524 138740
rect 484876 138740 484932 141708
rect 485100 139048 485156 142604
rect 485436 141764 485492 159628
rect 485884 158900 485940 160104
rect 485884 158834 485940 158844
rect 493948 157556 494004 160104
rect 493948 157490 494004 157500
rect 494732 160076 495208 160132
rect 495404 160076 495544 160132
rect 499688 160076 500612 160132
rect 500808 160076 501228 160132
rect 502124 160132 502180 160142
rect 493052 155652 493108 155662
rect 491372 155540 491428 155550
rect 485436 141698 485492 141708
rect 486332 152292 486388 152302
rect 486332 140420 486388 152236
rect 486332 139076 486388 140364
rect 491372 140308 491428 155484
rect 491372 139076 491428 140252
rect 485800 139020 486388 139076
rect 490952 139020 491428 139076
rect 491596 150612 491652 150622
rect 491596 140868 491652 150556
rect 491596 139076 491652 140812
rect 493052 140532 493108 155596
rect 493052 139076 493108 140476
rect 491596 139020 491960 139076
rect 492856 139020 493108 139076
rect 493388 147028 493444 147038
rect 493388 140756 493444 146972
rect 494732 141876 494788 160076
rect 494732 141810 494788 141820
rect 495404 142996 495460 160076
rect 493388 139048 493444 140700
rect 495404 139188 495460 142940
rect 496860 145796 496916 145806
rect 495516 142212 495572 142222
rect 495516 141876 495572 142156
rect 495516 141810 495572 141820
rect 495404 139122 495460 139132
rect 496860 139076 496916 145740
rect 500556 142884 500612 160076
rect 501228 160066 501284 160076
rect 500556 142818 500612 142828
rect 498988 142324 499044 142334
rect 498988 140196 499044 142268
rect 501452 142324 501508 160104
rect 502180 160076 502292 160132
rect 502600 160076 503972 160132
rect 504280 160076 505652 160132
rect 505960 160076 507332 160132
rect 502124 160066 502180 160076
rect 501452 142258 501508 142268
rect 498988 140130 499044 140140
rect 500668 141316 500724 141326
rect 500668 139188 500724 141260
rect 502236 141316 502292 160076
rect 502236 141250 502292 141260
rect 503916 141428 503972 160076
rect 505596 141540 505652 160076
rect 505596 141474 505652 141484
rect 506604 152068 506660 152078
rect 503916 140980 503972 141372
rect 503916 140914 503972 140924
rect 500668 139122 500724 139132
rect 506604 139048 506660 152012
rect 507276 141652 507332 160076
rect 512316 159572 512372 160104
rect 512316 159506 512372 159516
rect 520828 160076 522088 160132
rect 524188 160076 525560 160132
rect 520828 145796 520884 160076
rect 524188 147028 524244 160076
rect 526092 155652 526148 160104
rect 526092 155586 526148 155596
rect 526988 150612 527044 160104
rect 527996 155540 528052 160104
rect 527996 155474 528052 155484
rect 533148 152292 533204 160104
rect 533148 152226 533204 152236
rect 533372 160076 533848 160132
rect 526988 150546 527044 150556
rect 533372 149548 533428 160076
rect 534604 156212 534660 160104
rect 542892 157780 542948 160104
rect 542892 157714 542948 157724
rect 543004 160076 543480 160132
rect 543676 160076 543928 160132
rect 543004 156436 543060 160076
rect 534604 156146 534660 156156
rect 542556 156380 543060 156436
rect 542556 150500 542612 156380
rect 542556 150434 542612 150444
rect 543676 149548 543732 160076
rect 544348 152180 544404 160104
rect 544348 152114 544404 152124
rect 544572 160076 544824 160132
rect 524188 146962 524244 146972
rect 532588 149492 533428 149548
rect 542668 149492 543732 149548
rect 520828 145730 520884 145740
rect 532588 143892 532644 149492
rect 542668 145684 542724 149492
rect 544572 147140 544628 160076
rect 545468 157668 545524 160104
rect 545468 157602 545524 157612
rect 552076 159012 552132 159022
rect 544572 147074 544628 147084
rect 542668 145618 542724 145628
rect 532588 143826 532644 143836
rect 533036 145572 533092 145582
rect 524972 143780 525028 143790
rect 523404 142996 523460 143006
rect 519260 142884 519316 142894
rect 517468 142324 517524 142334
rect 507276 141586 507332 141596
rect 512988 141652 513044 141662
rect 512988 139048 513044 141596
rect 514668 141540 514724 141550
rect 514668 139048 514724 141484
rect 516348 141428 516404 141438
rect 516348 139048 516404 141372
rect 517468 139048 517524 142268
rect 518140 141316 518196 141326
rect 518140 139048 518196 141260
rect 519260 139048 519316 142828
rect 523404 139048 523460 142940
rect 523740 142212 523796 142222
rect 523740 139048 523796 142156
rect 524972 139048 525028 143724
rect 533036 139048 533092 145516
rect 535724 145460 535780 145470
rect 534156 142100 534212 142110
rect 533820 140644 533876 140654
rect 533820 139048 533876 140588
rect 534156 139048 534212 142044
rect 534940 141764 534996 141774
rect 534604 141204 534660 141214
rect 534604 139048 534660 141148
rect 534940 139048 534996 141708
rect 535724 139048 535780 145404
rect 543900 143668 543956 143678
rect 543900 139048 543956 143612
rect 545356 141988 545412 141998
rect 544684 141204 544740 141214
rect 544684 139048 544740 141148
rect 545356 139048 545412 141932
rect 496860 139010 496916 139020
rect 475244 138684 475496 138712
rect 475244 138628 475300 138684
rect 484876 138674 484932 138684
rect 475244 138562 475300 138572
rect 460236 36082 460292 36092
rect 460684 39508 460740 39518
rect 459452 4162 459508 4172
rect 460684 480 460740 39452
rect 489244 38052 489300 38062
rect 466396 6020 466452 6030
rect 466396 480 466452 5964
rect 472108 4676 472164 4686
rect 472108 480 472164 4620
rect 477820 4564 477876 4574
rect 477820 480 477876 4508
rect 483532 4452 483588 4462
rect 483532 480 483588 4396
rect 489244 480 489300 37996
rect 512092 37940 512148 37950
rect 506380 24388 506436 24398
rect 500668 5908 500724 5918
rect 494956 4340 495012 4350
rect 494956 480 495012 4284
rect 500668 480 500724 5852
rect 506380 480 506436 24332
rect 512092 480 512148 37884
rect 534940 37828 534996 37838
rect 517804 34468 517860 34478
rect 517804 480 517860 34412
rect 529228 32788 529284 32798
rect 523516 4228 523572 4238
rect 523516 480 523572 4172
rect 529228 480 529284 32732
rect 534940 480 534996 37772
rect 540652 36148 540708 36158
rect 540652 480 540708 36092
rect 546588 4228 546644 4238
rect 546588 480 546644 4172
rect 552076 480 552132 158956
rect 553532 157892 553588 160104
rect 553532 157826 553588 157836
rect 554428 156324 554484 160104
rect 554316 156268 554484 156324
rect 554316 150388 554372 156268
rect 555100 155428 555156 160104
rect 555100 155362 555156 155372
rect 554316 150322 554372 150332
rect 559468 4340 559524 379036
rect 590492 378868 590548 378878
rect 559468 4274 559524 4284
rect 559580 375508 559636 375518
rect 558012 4228 558068 4238
rect 558012 480 558068 4172
rect 559580 4228 559636 375452
rect 559580 4162 559636 4172
rect 563500 373828 563556 373838
rect 563500 480 563556 373772
rect 569212 372148 569268 372158
rect 565292 278292 565348 278302
rect 565292 7140 565348 278236
rect 568652 269668 568708 269678
rect 568652 139300 568708 269612
rect 568652 139234 568708 139244
rect 565292 7074 565348 7084
rect 569212 480 569268 372092
rect 574924 368900 574980 368910
rect 570332 276500 570388 276510
rect 570332 178948 570388 276444
rect 570332 178882 570388 178892
rect 574924 480 574980 368844
rect 590492 324548 590548 378812
rect 590604 364196 590660 380492
rect 590604 364130 590660 364140
rect 590492 324482 590548 324492
rect 590604 278180 590660 278190
rect 580636 273140 580692 273150
rect 580636 480 580692 273084
rect 582540 266420 582596 266430
rect 582540 480 582596 266364
rect 584444 264852 584500 264862
rect 584444 480 584500 264796
rect 590492 264628 590548 264638
rect 590492 47012 590548 264572
rect 590604 165956 590660 278124
rect 590716 268100 590772 268110
rect 590716 245252 590772 268044
rect 590716 245186 590772 245196
rect 590604 165890 590660 165900
rect 590604 160468 590660 160478
rect 590604 86660 590660 160412
rect 590604 86594 590660 86604
rect 590492 46946 590548 46956
rect 207452 392 207704 480
rect 209356 392 209608 480
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 392 211540 480
rect 211288 -960 211512 392
rect 213192 -960 213416 480
rect 215096 392 215348 480
rect 215096 -960 215320 392
rect 217000 -960 217224 480
rect 218904 -960 219128 480
rect 220808 392 221060 480
rect 220808 -960 221032 392
rect 222712 -960 222936 480
rect 224616 -960 224840 480
rect 226520 392 226772 480
rect 226520 -960 226744 392
rect 228424 -960 228648 480
rect 230328 -960 230552 480
rect 232232 392 232484 480
rect 232232 -960 232456 392
rect 234136 -960 234360 480
rect 236040 -960 236264 480
rect 237944 392 238196 480
rect 237944 -960 238168 392
rect 239848 -960 240072 480
rect 241752 -960 241976 480
rect 243656 392 243908 480
rect 243656 -960 243880 392
rect 245560 -960 245784 480
rect 247464 -960 247688 480
rect 249340 392 249592 480
rect 249368 -960 249592 392
rect 251272 -960 251496 480
rect 253176 -960 253400 480
rect 255052 392 255304 480
rect 255080 -960 255304 392
rect 256984 -960 257208 480
rect 258888 -960 259112 480
rect 260764 392 261016 480
rect 260792 -960 261016 392
rect 262696 -960 262920 480
rect 264600 -960 264824 480
rect 266504 392 266756 480
rect 266504 -960 266728 392
rect 268408 -960 268632 480
rect 270312 -960 270536 480
rect 272188 392 272440 480
rect 272216 -960 272440 392
rect 274120 -960 274344 480
rect 276024 -960 276248 480
rect 277900 392 278152 480
rect 277928 -960 278152 392
rect 279832 -960 280056 480
rect 281736 -960 281960 480
rect 283612 392 283864 480
rect 283640 -960 283864 392
rect 285544 -960 285768 480
rect 287448 -960 287672 480
rect 289324 392 289576 480
rect 289352 -960 289576 392
rect 291256 -960 291480 480
rect 293160 -960 293384 480
rect 295036 392 295288 480
rect 295064 -960 295288 392
rect 296968 -960 297192 480
rect 298872 -960 299096 480
rect 300748 392 301000 480
rect 300776 -960 301000 392
rect 302680 -960 302904 480
rect 304584 -960 304808 480
rect 306460 392 306712 480
rect 306488 -960 306712 392
rect 308392 -960 308616 480
rect 310296 -960 310520 480
rect 312172 392 312424 480
rect 312200 -960 312424 392
rect 314104 -960 314328 480
rect 316008 -960 316232 480
rect 317884 392 318136 480
rect 317912 -960 318136 392
rect 319816 -960 320040 480
rect 321720 -960 321944 480
rect 323596 392 323848 480
rect 323624 -960 323848 392
rect 325528 -960 325752 480
rect 327432 -960 327656 480
rect 329308 392 329560 480
rect 329336 -960 329560 392
rect 331240 -960 331464 480
rect 333144 -960 333368 480
rect 335048 392 335300 480
rect 335048 -960 335272 392
rect 336952 -960 337176 480
rect 338856 -960 339080 480
rect 340760 392 341012 480
rect 340760 -960 340984 392
rect 342664 -960 342888 480
rect 344568 -960 344792 480
rect 346472 392 346724 480
rect 346472 -960 346696 392
rect 348376 -960 348600 480
rect 350280 -960 350504 480
rect 352156 392 352408 480
rect 352184 -960 352408 392
rect 354088 -960 354312 480
rect 355992 -960 356216 480
rect 357868 392 358120 480
rect 357896 -960 358120 392
rect 359800 -960 360024 480
rect 361704 -960 361928 480
rect 363580 392 363832 480
rect 363608 -960 363832 392
rect 365512 -960 365736 480
rect 367416 -960 367640 480
rect 369292 392 369544 480
rect 369320 -960 369544 392
rect 371224 -960 371448 480
rect 373128 -960 373352 480
rect 375004 392 375256 480
rect 375032 -960 375256 392
rect 376936 -960 377160 480
rect 378840 -960 379064 480
rect 380716 392 380968 480
rect 380744 -960 380968 392
rect 382648 -960 382872 480
rect 384552 -960 384776 480
rect 386428 392 386680 480
rect 386456 -960 386680 392
rect 388360 -960 388584 480
rect 390264 -960 390488 480
rect 392140 392 392392 480
rect 392168 -960 392392 392
rect 394072 -960 394296 480
rect 395976 -960 396200 480
rect 397852 392 398104 480
rect 397880 -960 398104 392
rect 399784 -960 400008 480
rect 401688 -960 401912 480
rect 403564 392 403816 480
rect 403592 -960 403816 392
rect 405496 -960 405720 480
rect 407400 -960 407624 480
rect 409276 392 409528 480
rect 409304 -960 409528 392
rect 411208 -960 411432 480
rect 413112 -960 413336 480
rect 414988 392 415240 480
rect 415016 -960 415240 392
rect 416920 -960 417144 480
rect 418824 -960 419048 480
rect 420700 392 420952 480
rect 420728 -960 420952 392
rect 422632 -960 422856 480
rect 424536 -960 424760 480
rect 426412 392 426664 480
rect 426440 -960 426664 392
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432124 392 432376 480
rect 432152 -960 432376 392
rect 434056 -960 434280 480
rect 435960 -960 436184 480
rect 437836 392 438088 480
rect 437864 -960 438088 392
rect 439768 -960 439992 480
rect 441672 -960 441896 480
rect 443576 392 443828 480
rect 443576 -960 443800 392
rect 445480 -960 445704 480
rect 447384 -960 447608 480
rect 449260 392 449512 480
rect 449288 -960 449512 392
rect 451192 -960 451416 480
rect 453096 -960 453320 480
rect 454972 392 455224 480
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458808 -960 459032 480
rect 460684 392 460936 480
rect 460712 -960 460936 392
rect 462616 -960 462840 480
rect 464520 -960 464744 480
rect 466396 392 466648 480
rect 466424 -960 466648 392
rect 468328 -960 468552 480
rect 470232 -960 470456 480
rect 472108 392 472360 480
rect 472136 -960 472360 392
rect 474040 -960 474264 480
rect 475944 -960 476168 480
rect 477820 392 478072 480
rect 477848 -960 478072 392
rect 479752 -960 479976 480
rect 481656 -960 481880 480
rect 483532 392 483784 480
rect 483560 -960 483784 392
rect 485464 -960 485688 480
rect 487368 -960 487592 480
rect 489244 392 489496 480
rect 489272 -960 489496 392
rect 491176 -960 491400 480
rect 493080 -960 493304 480
rect 494956 392 495208 480
rect 494984 -960 495208 392
rect 496888 -960 497112 480
rect 498792 -960 499016 480
rect 500668 392 500920 480
rect 500696 -960 500920 392
rect 502600 -960 502824 480
rect 504504 -960 504728 480
rect 506380 392 506632 480
rect 506408 -960 506632 392
rect 508312 -960 508536 480
rect 510216 -960 510440 480
rect 512092 392 512344 480
rect 512120 -960 512344 392
rect 514024 -960 514248 480
rect 515928 -960 516152 480
rect 517804 392 518056 480
rect 517832 -960 518056 392
rect 519736 -960 519960 480
rect 521640 -960 521864 480
rect 523516 392 523768 480
rect 523544 -960 523768 392
rect 525448 -960 525672 480
rect 527352 -960 527576 480
rect 529228 392 529480 480
rect 529256 -960 529480 392
rect 531160 -960 531384 480
rect 533064 -960 533288 480
rect 534940 392 535192 480
rect 534968 -960 535192 392
rect 536872 -960 537096 480
rect 538776 -960 539000 480
rect 540652 392 540904 480
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544488 -960 544712 480
rect 546392 392 546644 480
rect 546392 -960 546616 392
rect 548296 -960 548520 480
rect 550200 -960 550424 480
rect 552076 392 552328 480
rect 552104 -960 552328 392
rect 554008 -960 554232 480
rect 555912 -960 556136 480
rect 557816 392 558068 480
rect 557816 -960 558040 392
rect 559720 -960 559944 480
rect 561624 -960 561848 480
rect 563500 392 563752 480
rect 563528 -960 563752 392
rect 565432 -960 565656 480
rect 567336 -960 567560 480
rect 569212 392 569464 480
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573048 -960 573272 480
rect 574924 392 575176 480
rect 574952 -960 575176 392
rect 576856 -960 577080 480
rect 578760 -960 578984 480
rect 580636 392 580888 480
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 55356 590604 55412 590660
rect 33292 590492 33348 590548
rect 11004 563612 11060 563668
rect 50316 588812 50372 588868
rect 4284 516572 4340 516628
rect 4172 502460 4228 502516
rect 20972 486332 21028 486388
rect 15932 466172 15988 466228
rect 14252 464492 14308 464548
rect 4284 452732 4340 452788
rect 4396 460124 4452 460180
rect 12572 457772 12628 457828
rect 7532 449372 7588 449428
rect 4396 436156 4452 436212
rect 4956 446012 5012 446068
rect 4956 436044 5012 436100
rect 4172 435932 4228 435988
rect 4620 429772 4676 429828
rect 4396 429660 4452 429716
rect 4172 429548 4228 429604
rect 4620 418012 4676 418068
rect 4396 389676 4452 389732
rect 4172 375676 4228 375732
rect 4284 271516 4340 271572
rect 4172 269724 4228 269780
rect 4508 266252 4564 266308
rect 4396 264684 4452 264740
rect 4508 220444 4564 220500
rect 4396 192220 4452 192276
rect 4284 177996 4340 178052
rect 4172 163996 4228 164052
rect 4172 160636 4228 160692
rect 4172 135772 4228 135828
rect 7532 65212 7588 65268
rect 11340 141932 11396 141988
rect 12572 93212 12628 93268
rect 14252 50876 14308 50932
rect 19292 446012 19348 446068
rect 15932 8540 15988 8596
rect 17612 211036 17668 211092
rect 15372 4396 15428 4452
rect 13356 4284 13412 4340
rect 19292 107324 19348 107380
rect 20972 36764 21028 36820
rect 22652 467852 22708 467908
rect 17612 4284 17668 4340
rect 18956 24332 19012 24388
rect 17276 4172 17332 4228
rect 50204 420364 50260 420420
rect 48636 416332 48692 416388
rect 48412 401548 48468 401604
rect 26012 286748 26068 286804
rect 22652 22652 22708 22708
rect 24332 230972 24388 231028
rect 20860 13356 20916 13412
rect 24332 4172 24388 4228
rect 24668 217644 24724 217700
rect 22988 4060 23044 4116
rect 26012 24332 26068 24388
rect 27692 286636 27748 286692
rect 27692 13356 27748 13412
rect 29372 285068 29428 285124
rect 32732 278348 32788 278404
rect 31052 214284 31108 214340
rect 29372 4284 29428 4340
rect 30604 4844 30660 4900
rect 26796 4172 26852 4228
rect 48412 257852 48468 257908
rect 48524 397516 48580 397572
rect 45612 254492 45668 254548
rect 32732 4844 32788 4900
rect 34412 252812 34468 252868
rect 31052 4060 31108 4116
rect 32508 4284 32564 4340
rect 42812 251132 42868 251188
rect 37996 224252 38052 224308
rect 34412 4284 34468 4340
rect 34524 4508 34580 4564
rect 40124 4844 40180 4900
rect 42028 4284 42084 4340
rect 44492 232652 44548 232708
rect 44492 4844 44548 4900
rect 42812 4284 42868 4340
rect 48524 222684 48580 222740
rect 47852 219212 47908 219268
rect 49980 414988 50036 415044
rect 49980 284956 50036 285012
rect 50092 402892 50148 402948
rect 50092 266364 50148 266420
rect 49532 246092 49588 246148
rect 48636 215852 48692 215908
rect 49420 222572 49476 222628
rect 47852 4284 47908 4340
rect 47740 4172 47796 4228
rect 55356 583772 55412 583828
rect 53676 582092 53732 582148
rect 51884 578732 51940 578788
rect 50316 342412 50372 342468
rect 51772 398860 51828 398916
rect 51884 314188 51940 314244
rect 51996 432124 52052 432180
rect 51772 283276 51828 283332
rect 50204 227612 50260 227668
rect 51212 234332 51268 234388
rect 53676 339724 53732 339780
rect 55244 430332 55300 430388
rect 53676 324268 53732 324324
rect 51996 160412 52052 160468
rect 53228 229292 53284 229348
rect 51212 4508 51268 4564
rect 49532 4172 49588 4228
rect 58716 582204 58772 582260
rect 58492 572124 58548 572180
rect 57036 566972 57092 567028
rect 56924 430108 56980 430164
rect 56812 427308 56868 427364
rect 56700 427196 56756 427252
rect 56700 410956 56756 411012
rect 56812 409612 56868 409668
rect 56924 405580 56980 405636
rect 56924 400204 56980 400260
rect 56700 396172 56756 396228
rect 55356 341068 55412 341124
rect 56252 394828 56308 394884
rect 56700 354396 56756 354452
rect 56812 393484 56868 393540
rect 56252 324268 56308 324324
rect 56812 307356 56868 307412
rect 55244 212828 55300 212884
rect 55356 300748 55412 300804
rect 53676 212604 53732 212660
rect 56700 300748 56756 300804
rect 58380 423052 58436 423108
rect 58268 419020 58324 419076
rect 57036 318220 57092 318276
rect 58156 417676 58212 417732
rect 56924 300076 56980 300132
rect 56700 291788 56756 291844
rect 56812 299404 56868 299460
rect 57036 298060 57092 298116
rect 56812 276444 56868 276500
rect 56924 294028 56980 294084
rect 55356 33628 55412 33684
rect 56252 273084 56308 273140
rect 55356 4956 55412 5012
rect 56924 269836 56980 269892
rect 58156 288092 58212 288148
rect 58268 284844 58324 284900
rect 57036 269612 57092 269668
rect 58492 343756 58548 343812
rect 58604 565404 58660 565460
rect 58604 316876 58660 316932
rect 99484 590716 99540 590772
rect 121324 570332 121380 570388
rect 121772 572012 121828 572068
rect 77308 565292 77364 565348
rect 104412 488012 104468 488068
rect 101724 437612 101780 437668
rect 99036 434252 99092 434308
rect 90972 432908 91028 432964
rect 66780 432124 66836 432180
rect 64092 432012 64148 432068
rect 60396 431900 60452 431956
rect 60060 425068 60116 425124
rect 58716 315532 58772 315588
rect 59612 354396 59668 354452
rect 58380 217532 58436 217588
rect 58716 286524 58772 286580
rect 58604 214172 58660 214228
rect 56252 4956 56308 5012
rect 57148 139356 57204 139412
rect 59836 307356 59892 307412
rect 59612 212716 59668 212772
rect 59724 286412 59780 286468
rect 58716 37884 58772 37940
rect 58940 211148 58996 211204
rect 58604 3948 58660 4004
rect 60172 423836 60228 423892
rect 60172 284732 60228 284788
rect 60284 421596 60340 421652
rect 60284 283164 60340 283220
rect 60060 283052 60116 283108
rect 88284 432012 88340 432068
rect 72156 431900 72212 431956
rect 69468 430220 69524 430276
rect 82908 431900 82964 431956
rect 77532 431788 77588 431844
rect 85596 431900 85652 431956
rect 96348 432572 96404 432628
rect 93660 430220 93716 430276
rect 109788 484652 109844 484708
rect 107100 432684 107156 432740
rect 120540 469532 120596 469588
rect 117852 433468 117908 433524
rect 112476 432236 112532 432292
rect 115164 432124 115220 432180
rect 165676 590828 165732 590884
rect 143388 555212 143444 555268
rect 153692 557788 153748 557844
rect 144732 500668 144788 500724
rect 136668 499772 136724 499828
rect 133980 498092 134036 498148
rect 131292 437724 131348 437780
rect 121772 432684 121828 432740
rect 123228 433580 123284 433636
rect 128604 432348 128660 432404
rect 142044 434476 142100 434532
rect 139356 434364 139412 434420
rect 150108 498204 150164 498260
rect 147420 494732 147476 494788
rect 173740 557788 173796 557844
rect 231756 591052 231812 591108
rect 209804 590940 209860 590996
rect 320124 591276 320180 591332
rect 298060 591164 298116 591220
rect 279692 590940 279748 590996
rect 275996 590156 276052 590212
rect 278012 590156 278068 590212
rect 253932 588924 253988 588980
rect 187516 555324 187572 555380
rect 274652 554428 274708 554484
rect 201292 554316 201348 554372
rect 216748 551516 216804 551572
rect 215740 548828 215796 548884
rect 215180 543452 215236 543508
rect 214508 510748 214564 510804
rect 214396 505708 214452 505764
rect 160860 501452 160916 501508
rect 153692 476252 153748 476308
rect 155484 499884 155540 499940
rect 152796 444332 152852 444388
rect 158172 437836 158228 437892
rect 176988 500556 177044 500612
rect 162764 486332 162820 486388
rect 167244 446012 167300 446068
rect 171500 499996 171556 500052
rect 163548 433356 163604 433412
rect 166236 433356 166292 433412
rect 169596 433356 169652 433412
rect 176204 467852 176260 467908
rect 171724 449372 171780 449428
rect 174300 449372 174356 449428
rect 179676 493052 179732 493108
rect 180684 457772 180740 457828
rect 182364 491372 182420 491428
rect 198604 496524 198660 496580
rect 202412 497196 202468 497252
rect 194124 496412 194180 496468
rect 189644 466172 189700 466228
rect 185164 464492 185220 464548
rect 187740 451052 187796 451108
rect 185052 437948 185108 438004
rect 212044 469532 212100 469588
rect 207564 452844 207620 452900
rect 202412 444332 202468 444388
rect 190428 439292 190484 439348
rect 214396 437836 214452 437892
rect 215068 508508 215124 508564
rect 214844 502796 214900 502852
rect 215068 501452 215124 501508
rect 214844 499884 214900 499940
rect 215292 540764 215348 540820
rect 215404 538076 215460 538132
rect 215404 501676 215460 501732
rect 215516 516572 215572 516628
rect 215516 499772 215572 499828
rect 215628 513884 215684 513940
rect 215628 513212 215684 513268
rect 215628 498092 215684 498148
rect 215292 493052 215348 493108
rect 215180 491372 215236 491428
rect 215740 451052 215796 451108
rect 217532 550172 217588 550228
rect 217308 532700 217364 532756
rect 217084 530012 217140 530068
rect 216748 439292 216804 439348
rect 216860 521612 216916 521668
rect 214508 437724 214564 437780
rect 216860 434476 216916 434532
rect 216972 519932 217028 519988
rect 217084 498204 217140 498260
rect 217196 527436 217252 527492
rect 217308 501564 217364 501620
rect 217756 549388 217812 549444
rect 217756 527436 217812 527492
rect 218428 546140 218484 546196
rect 217532 524636 217588 524692
rect 217532 500668 217588 500724
rect 217196 494732 217252 494788
rect 218540 535388 218596 535444
rect 218540 449372 218596 449428
rect 246876 452844 246932 452900
rect 218428 437948 218484 438004
rect 216972 434364 217028 434420
rect 209244 432572 209300 432628
rect 206556 432460 206612 432516
rect 203868 430556 203924 430612
rect 193116 430332 193172 430388
rect 201180 430332 201236 430388
rect 244188 430780 244244 430836
rect 219996 430668 220052 430724
rect 214620 430444 214676 430500
rect 212828 429996 212884 430052
rect 265692 433356 265748 433412
rect 257628 431004 257684 431060
rect 254940 430892 254996 430948
rect 268716 433356 268772 433412
rect 272636 432684 272692 432740
rect 80220 429436 80276 429492
rect 74844 429324 74900 429380
rect 125916 429212 125972 429268
rect 217308 429212 217364 429268
rect 249564 429212 249620 429268
rect 252252 429212 252308 429268
rect 260316 429212 260372 429268
rect 263004 429212 263060 429268
rect 60620 428540 60676 428596
rect 270620 422380 270676 422436
rect 269500 409948 269556 410004
rect 269388 405692 269444 405748
rect 60396 278124 60452 278180
rect 60620 300076 60676 300132
rect 59836 212940 59892 212996
rect 63756 290108 63812 290164
rect 60620 212492 60676 212548
rect 61180 286860 61236 286916
rect 60284 210924 60340 210980
rect 60172 210812 60228 210868
rect 59724 37772 59780 37828
rect 59948 209468 60004 209524
rect 59948 4284 60004 4340
rect 60060 209356 60116 209412
rect 60172 4396 60228 4452
rect 67228 285068 67284 285124
rect 71260 286748 71316 286804
rect 73276 286636 73332 286692
rect 69244 230972 69300 231028
rect 81340 278348 81396 278404
rect 83356 252812 83412 252868
rect 85372 234332 85428 234388
rect 89404 232652 89460 232708
rect 91196 283276 91252 283332
rect 87388 224252 87444 224308
rect 79324 219212 79380 219268
rect 87164 222684 87220 222740
rect 77308 217644 77364 217700
rect 75292 214284 75348 214340
rect 65212 211036 65268 211092
rect 66668 213276 66724 213332
rect 62972 209916 63028 209972
rect 75068 212940 75124 212996
rect 71036 212828 71092 212884
rect 83132 212716 83188 212772
rect 79100 212604 79156 212660
rect 93436 254492 93492 254548
rect 91420 251132 91476 251188
rect 95452 246092 95508 246148
rect 96572 285628 96628 285684
rect 97468 285628 97524 285684
rect 96572 222572 96628 222628
rect 99260 257852 99316 257908
rect 95228 212492 95284 212548
rect 103516 286860 103572 286916
rect 101500 273084 101556 273140
rect 99484 229292 99540 229348
rect 103292 266364 103348 266420
rect 105532 211148 105588 211204
rect 107324 284956 107380 285012
rect 107548 209468 107604 209524
rect 111356 215852 111412 215908
rect 111580 210924 111636 210980
rect 113596 210812 113652 210868
rect 115388 288092 115444 288148
rect 115612 281372 115668 281428
rect 119644 286524 119700 286580
rect 117628 227724 117684 227780
rect 119420 284844 119476 284900
rect 123676 286412 123732 286468
rect 127708 286300 127764 286356
rect 125692 285628 125748 285684
rect 127484 283164 127540 283220
rect 121660 214172 121716 214228
rect 123452 227612 123508 227668
rect 131740 286524 131796 286580
rect 129724 257964 129780 258020
rect 135772 286300 135828 286356
rect 137788 286188 137844 286244
rect 139804 285628 139860 285684
rect 143836 286524 143892 286580
rect 147868 286188 147924 286244
rect 145852 285964 145908 286020
rect 149884 285740 149940 285796
rect 141820 285628 141876 285684
rect 153916 285628 153972 285684
rect 155932 285628 155988 285684
rect 157052 285628 157108 285684
rect 151900 285068 151956 285124
rect 151676 284844 151732 284900
rect 133756 231084 133812 231140
rect 135548 284732 135604 284788
rect 131516 217532 131572 217588
rect 143612 284732 143668 284788
rect 139580 283052 139636 283108
rect 147644 283052 147700 283108
rect 157948 285628 158004 285684
rect 159740 285628 159796 285684
rect 157052 222572 157108 222628
rect 155708 217532 155764 217588
rect 159740 212492 159796 212548
rect 109564 209356 109620 209412
rect 166012 285628 166068 285684
rect 163996 283276 164052 283332
rect 167804 266364 167860 266420
rect 163772 222572 163828 222628
rect 170044 286860 170100 286916
rect 174076 285628 174132 285684
rect 176092 285628 176148 285684
rect 178108 285628 178164 285684
rect 180124 230972 180180 231028
rect 179900 212828 179956 212884
rect 172060 212716 172116 212772
rect 175868 212716 175924 212772
rect 168028 210812 168084 210868
rect 171836 212604 171892 212660
rect 184156 285628 184212 285684
rect 186172 285628 186228 285684
rect 190204 286412 190260 286468
rect 188188 285628 188244 285684
rect 194236 286636 194292 286692
rect 191548 285628 191604 285684
rect 196252 285628 196308 285684
rect 200284 286972 200340 287028
rect 202300 285740 202356 285796
rect 198268 285628 198324 285684
rect 206332 286748 206388 286804
rect 204316 285628 204372 285684
rect 210364 286860 210420 286916
rect 212380 286524 212436 286580
rect 208348 285628 208404 285684
rect 214396 285628 214452 285684
rect 216412 285628 216468 285684
rect 220444 286412 220500 286468
rect 218428 285628 218484 285684
rect 221788 285628 221844 285684
rect 196028 284956 196084 285012
rect 191996 283164 192052 283220
rect 187964 224252 188020 224308
rect 182140 210924 182196 210980
rect 183932 214172 183988 214228
rect 200060 283276 200116 283332
rect 226492 285628 226548 285684
rect 230524 285740 230580 285796
rect 228508 285628 228564 285684
rect 231868 285628 231924 285684
rect 224476 281372 224532 281428
rect 228284 261324 228340 261380
rect 222572 260428 222628 260484
rect 216188 259644 216244 259700
rect 208124 258748 208180 258804
rect 204092 257852 204148 257908
rect 212156 215852 212212 215908
rect 220220 213276 220276 213332
rect 222572 213276 222628 213332
rect 224252 259756 224308 259812
rect 232316 258860 232372 258916
rect 236572 286412 236628 286468
rect 238588 285628 238644 285684
rect 240604 285628 240660 285684
rect 244636 285740 244692 285796
rect 242620 285628 242676 285684
rect 246876 285628 246932 285684
rect 250684 286300 250740 286356
rect 249228 285628 249284 285684
rect 254716 286412 254772 286468
rect 252140 285628 252196 285684
rect 256732 285628 256788 285684
rect 258748 285628 258804 285684
rect 262780 285852 262836 285908
rect 264796 285740 264852 285796
rect 260428 285628 260484 285684
rect 266812 285628 266868 285684
rect 248444 269948 248500 270004
rect 234556 210812 234612 210868
rect 236348 261436 236404 261492
rect 240380 254492 240436 254548
rect 244412 217644 244468 217700
rect 264572 268156 264628 268212
rect 260540 222684 260596 222740
rect 256508 215964 256564 216020
rect 252476 214284 252532 214340
rect 268604 266476 268660 266532
rect 270508 408940 270564 408996
rect 269500 266364 269556 266420
rect 269612 347788 269668 347844
rect 269388 217532 269444 217588
rect 269836 306236 269892 306292
rect 269724 303996 269780 304052
rect 269724 289772 269780 289828
rect 270732 421036 270788 421092
rect 270844 419692 270900 419748
rect 272188 414316 272244 414372
rect 270844 284956 270900 285012
rect 270956 404908 271012 404964
rect 270956 284844 271012 284900
rect 271292 334348 271348 334404
rect 270732 283276 270788 283332
rect 270620 257852 270676 257908
rect 270508 222572 270564 222628
rect 269836 212716 269892 212772
rect 272300 412972 272356 413028
rect 272412 411628 272468 411684
rect 272524 407596 272580 407652
rect 272972 432572 273028 432628
rect 273980 418348 274036 418404
rect 272972 397292 273028 397348
rect 273868 415660 273924 415716
rect 272636 388780 272692 388836
rect 272972 381388 273028 381444
rect 272972 369964 273028 370020
rect 272524 347788 272580 347844
rect 272412 334348 272468 334404
rect 273084 335020 273140 335076
rect 272300 306236 272356 306292
rect 272972 333676 273028 333732
rect 272300 302764 272356 302820
rect 272300 291452 272356 291508
rect 273084 279692 273140 279748
rect 273196 332332 273252 332388
rect 273196 276556 273252 276612
rect 273308 328300 273364 328356
rect 273532 326956 273588 327012
rect 273420 325612 273476 325668
rect 273756 318892 273812 318948
rect 273756 279916 273812 279972
rect 273532 279804 273588 279860
rect 273420 278348 273476 278404
rect 273308 273196 273364 273252
rect 272972 257852 273028 257908
rect 274092 402220 274148 402276
rect 274652 398188 274708 398244
rect 274764 432460 274820 432516
rect 274764 383852 274820 383908
rect 275548 417004 275604 417060
rect 274092 284732 274148 284788
rect 273980 283164 274036 283220
rect 275660 403564 275716 403620
rect 278124 553532 278180 553588
rect 278124 400876 278180 400932
rect 299964 590940 300020 590996
rect 298284 590380 298340 590436
rect 279804 562156 279860 562212
rect 291452 553420 291508 553476
rect 289772 552860 289828 552916
rect 279804 434252 279860 434308
rect 284732 496524 284788 496580
rect 279692 381836 279748 381892
rect 279804 431900 279860 431956
rect 288092 496412 288148 496468
rect 284732 402892 284788 402948
rect 284844 432236 284900 432292
rect 279804 380492 279860 380548
rect 278012 380156 278068 380212
rect 288092 402780 288148 402836
rect 296492 549724 296548 549780
rect 291452 399532 291508 399588
rect 293132 549612 293188 549668
rect 293132 396844 293188 396900
rect 294812 549276 294868 549332
rect 294812 394156 294868 394212
rect 294924 474236 294980 474292
rect 289772 390124 289828 390180
rect 284844 379596 284900 379652
rect 295036 433580 295092 433636
rect 295260 433468 295316 433524
rect 295148 432124 295204 432180
rect 295148 401436 295204 401492
rect 295260 399756 295316 399812
rect 295036 398076 295092 398132
rect 298172 548716 298228 548772
rect 298060 429772 298116 429828
rect 298060 401324 298116 401380
rect 296492 392812 296548 392868
rect 299852 551068 299908 551124
rect 298284 484652 298340 484708
rect 298396 488348 298452 488404
rect 298172 391468 298228 391524
rect 298284 432348 298340 432404
rect 298844 436044 298900 436100
rect 298620 435932 298676 435988
rect 298396 401212 298452 401268
rect 298508 429660 298564 429716
rect 298620 402556 298676 402612
rect 298844 402220 298900 402276
rect 341964 572124 342020 572180
rect 386092 590380 386148 590436
rect 408268 588812 408324 588868
rect 364028 566972 364084 567028
rect 451276 591164 451332 591220
rect 430220 565404 430276 565460
rect 449372 591052 449428 591108
rect 416780 554428 416836 554484
rect 318220 553308 318276 553364
rect 313292 553196 313348 553252
rect 303436 553084 303492 553140
rect 308364 552972 308420 553028
rect 382396 551516 382452 551572
rect 377356 551404 377412 551460
rect 372428 551292 372484 551348
rect 367500 551180 367556 551236
rect 367164 549948 367220 550004
rect 372428 549836 372484 549892
rect 377356 550172 377412 550228
rect 362572 549500 362628 549556
rect 323148 549388 323204 549444
rect 328076 549388 328132 549444
rect 333004 549388 333060 549444
rect 337932 549388 337988 549444
rect 342860 549388 342916 549444
rect 347788 549388 347844 549444
rect 352716 549388 352772 549444
rect 357644 549388 357700 549444
rect 406924 551068 406980 551124
rect 397068 549836 397124 549892
rect 426636 553532 426692 553588
rect 421708 553420 421764 553476
rect 436492 552860 436548 552916
rect 430780 550060 430836 550116
rect 387212 549724 387268 549780
rect 392812 549724 392868 549780
rect 382284 549388 382340 549444
rect 392140 549388 392196 549444
rect 411852 549612 411908 549668
rect 392812 549388 392868 549444
rect 401996 549276 402052 549332
rect 431340 549276 431396 549332
rect 441420 549276 441476 549332
rect 301084 549052 301140 549108
rect 300972 548604 301028 548660
rect 300972 530012 301028 530068
rect 301084 508172 301140 508228
rect 299964 488012 300020 488068
rect 451052 590492 451108 590548
rect 449372 434364 449428 434420
rect 449484 553084 449540 553140
rect 301084 430780 301140 430836
rect 300860 427644 300916 427700
rect 300860 401100 300916 401156
rect 449708 449372 449764 449428
rect 451052 446124 451108 446180
rect 451164 553196 451220 553252
rect 464492 591276 464548 591332
rect 456204 590828 456260 590884
rect 456092 587132 456148 587188
rect 452284 572012 452340 572068
rect 452732 573020 452788 573076
rect 451276 449484 451332 449540
rect 451164 437612 451220 437668
rect 454412 563612 454468 563668
rect 452844 553308 452900 553364
rect 452844 446012 452900 446068
rect 452732 434252 452788 434308
rect 449484 429548 449540 429604
rect 301084 400428 301140 400484
rect 299852 395500 299908 395556
rect 298508 380268 298564 380324
rect 298284 380044 298340 380100
rect 294924 379484 294980 379540
rect 299068 378924 299124 378980
rect 454524 552972 454580 553028
rect 454524 439292 454580 439348
rect 456204 444332 456260 444388
rect 457772 590716 457828 590772
rect 456092 437836 456148 437892
rect 459564 590604 459620 590660
rect 459452 549276 459508 549332
rect 462812 588924 462868 588980
rect 461244 570332 461300 570388
rect 459564 449596 459620 449652
rect 461132 565292 461188 565348
rect 459452 448476 459508 448532
rect 457772 437724 457828 437780
rect 454412 377580 454468 377636
rect 456092 429996 456148 430052
rect 299068 376684 299124 376740
rect 294924 375340 294980 375396
rect 289772 373996 289828 374052
rect 284732 330988 284788 331044
rect 279020 309484 279076 309540
rect 278908 306796 278964 306852
rect 278796 305452 278852 305508
rect 275660 283052 275716 283108
rect 277676 300076 277732 300132
rect 275548 224252 275604 224308
rect 276668 264908 276724 264964
rect 273868 214172 273924 214228
rect 271516 212828 271572 212884
rect 271292 212604 271348 212660
rect 269612 212492 269668 212548
rect 272636 212492 272692 212548
rect 161980 209356 162036 209412
rect 69020 157724 69076 157780
rect 71708 157052 71764 157108
rect 73836 157724 73892 157780
rect 66332 156492 66388 156548
rect 70476 156492 70532 156548
rect 63868 155484 63924 155540
rect 74396 157164 74452 157220
rect 73836 155372 73892 155428
rect 70476 152124 70532 152180
rect 65436 150332 65492 150388
rect 64428 142268 64484 142324
rect 61180 139356 61236 139412
rect 63756 141148 63812 141204
rect 77084 148652 77140 148708
rect 76076 146972 76132 147028
rect 73500 145404 73556 145460
rect 74620 142156 74676 142212
rect 74172 141932 74228 141988
rect 75068 142044 75124 142100
rect 75516 141260 75572 141316
rect 82460 142156 82516 142212
rect 84252 143612 84308 143668
rect 79772 142044 79828 142100
rect 84924 142268 84980 142324
rect 85036 148652 85092 148708
rect 93212 155708 93268 155764
rect 90524 145516 90580 145572
rect 87836 143724 87892 143780
rect 90972 141708 91028 141764
rect 85036 141036 85092 141092
rect 85820 141372 85876 141428
rect 96908 155484 96964 155540
rect 95900 141708 95956 141764
rect 96460 141708 96516 141764
rect 91980 141484 92036 141540
rect 92764 141148 92820 141204
rect 93324 140588 93380 140644
rect 96460 140252 96516 140308
rect 97692 141484 97748 141540
rect 98588 141484 98644 141540
rect 100828 141148 100884 141204
rect 103964 140588 104020 140644
rect 106652 155596 106708 155652
rect 100828 140476 100884 140532
rect 97692 140364 97748 140420
rect 96908 139244 96964 139300
rect 112028 155484 112084 155540
rect 109340 148652 109396 148708
rect 106764 147084 106820 147140
rect 112588 143724 112644 143780
rect 117404 157276 117460 157332
rect 114716 143724 114772 143780
rect 116732 155708 116788 155764
rect 112588 142492 112644 142548
rect 114716 141148 114772 141204
rect 118188 148652 118244 148708
rect 116732 139804 116788 139860
rect 117516 147084 117572 147140
rect 117516 140812 117572 140868
rect 120092 147868 120148 147924
rect 123564 157164 123620 157220
rect 122668 141372 122724 141428
rect 119308 141148 119364 141204
rect 123340 147868 123396 147924
rect 123340 139020 123396 139076
rect 123564 141484 123620 141540
rect 125020 145628 125076 145684
rect 124348 141260 124404 141316
rect 124348 140700 124404 140756
rect 128156 141932 128212 141988
rect 129276 142604 129332 142660
rect 133532 155596 133588 155652
rect 133756 157276 133812 157332
rect 130956 142268 131012 142324
rect 133084 144060 133140 144116
rect 129276 141932 129332 141988
rect 125468 140700 125524 140756
rect 133756 139580 133812 139636
rect 133980 157052 134036 157108
rect 133980 141372 134036 141428
rect 134652 155372 134708 155428
rect 138908 155708 138964 155764
rect 141596 155372 141652 155428
rect 146972 159516 147028 159572
rect 149100 157276 149156 157332
rect 144284 152012 144340 152068
rect 146972 157164 147028 157220
rect 136220 145516 136276 145572
rect 146972 145404 147028 145460
rect 148428 148652 148484 148708
rect 143836 144396 143892 144452
rect 134652 141820 134708 141876
rect 134988 143724 135044 143780
rect 135660 143724 135716 143780
rect 144732 142716 144788 142772
rect 145404 142380 145460 142436
rect 145404 141148 145460 141204
rect 122668 138796 122724 138852
rect 118188 138684 118244 138740
rect 135436 138572 135492 138628
rect 142828 40236 142884 40292
rect 97020 39452 97076 39508
rect 72268 37884 72324 37940
rect 66556 4396 66612 4452
rect 60284 4172 60340 4228
rect 60844 4284 60900 4340
rect 60060 4060 60116 4116
rect 64652 4172 64708 4228
rect 62748 4060 62804 4116
rect 68684 4284 68740 4340
rect 70364 4172 70420 4228
rect 76076 37772 76132 37828
rect 74172 4060 74228 4116
rect 95116 36092 95172 36148
rect 83692 26012 83748 26068
rect 78204 4172 78260 4228
rect 80108 4172 80164 4228
rect 82012 4172 82068 4228
rect 87500 24332 87556 24388
rect 85820 4284 85876 4340
rect 91308 15932 91364 15988
rect 89628 5964 89684 6020
rect 93436 7532 93492 7588
rect 106540 37884 106596 37940
rect 104636 12572 104692 12628
rect 99036 7644 99092 7700
rect 101052 5852 101108 5908
rect 102956 4172 103012 4228
rect 110348 37772 110404 37828
rect 108668 4172 108724 4228
rect 119868 36204 119924 36260
rect 112476 4172 112532 4228
rect 114380 4172 114436 4228
rect 118188 4172 118244 4228
rect 116284 4060 116340 4116
rect 139132 5068 139188 5124
rect 133420 4732 133476 4788
rect 121996 4620 122052 4676
rect 127596 4508 127652 4564
rect 125804 4396 125860 4452
rect 123900 4284 123956 4340
rect 131516 4060 131572 4116
rect 129612 3948 129668 4004
rect 135324 4620 135380 4676
rect 137228 3388 137284 3444
rect 141036 4844 141092 4900
rect 146748 4956 146804 5012
rect 144844 4732 144900 4788
rect 148652 143948 148708 144004
rect 148876 143836 148932 143892
rect 149660 144396 149716 144452
rect 150332 147196 150388 147252
rect 149100 143612 149156 143668
rect 148876 4508 148932 4564
rect 148652 4284 148708 4340
rect 150444 145740 150500 145796
rect 152012 145404 152068 145460
rect 153692 156268 153748 156324
rect 157276 158844 157332 158900
rect 155036 156268 155092 156324
rect 155372 157052 155428 157108
rect 153692 144060 153748 144116
rect 154140 144172 154196 144228
rect 152348 143724 152404 143780
rect 152572 143724 152628 143780
rect 152012 4732 152068 4788
rect 150444 4396 150500 4452
rect 152460 4284 152516 4340
rect 152572 4060 152628 4116
rect 157276 4844 157332 4900
rect 157500 147084 157556 147140
rect 155372 4620 155428 4676
rect 160412 157276 160468 157332
rect 162092 156268 162148 156324
rect 160860 152348 160916 152404
rect 157724 145628 157780 145684
rect 159852 145628 159908 145684
rect 157500 4508 157556 4564
rect 157948 143612 158004 143668
rect 156156 4172 156212 4228
rect 165788 157164 165844 157220
rect 163100 156268 163156 156324
rect 168476 150332 168532 150388
rect 162092 146972 162148 147028
rect 174748 150444 174804 150500
rect 176092 152796 176148 152852
rect 171164 146972 171220 147028
rect 173516 145628 173572 145684
rect 165340 144060 165396 144116
rect 163772 142268 163828 142324
rect 164556 142268 164612 142324
rect 164556 141932 164612 141988
rect 164444 141260 164500 141316
rect 174188 142604 174244 142660
rect 174188 139692 174244 139748
rect 174636 142156 174692 142212
rect 174636 141596 174692 141652
rect 174972 142044 175028 142100
rect 175420 140700 175476 140756
rect 175420 139020 175476 139076
rect 179228 157276 179284 157332
rect 184604 152796 184660 152852
rect 181916 147868 181972 147924
rect 184268 147868 184324 147924
rect 176540 147084 176596 147140
rect 176316 142044 176372 142100
rect 176316 141708 176372 141764
rect 187292 145628 187348 145684
rect 188972 156268 189028 156324
rect 195356 157164 195412 157220
rect 192668 157052 192724 157108
rect 189980 156268 190036 156324
rect 200732 155820 200788 155876
rect 203420 152236 203476 152292
rect 198268 150556 198324 150612
rect 188972 144060 189028 144116
rect 208796 157388 208852 157444
rect 216860 157500 216916 157556
rect 214172 155484 214228 155540
rect 222236 152124 222292 152180
rect 222572 157276 222628 157332
rect 219548 150332 219604 150388
rect 211484 147308 211540 147364
rect 206108 144060 206164 144116
rect 206556 145516 206612 145572
rect 186396 142044 186452 142100
rect 185052 141148 185108 141204
rect 186396 141148 186452 141204
rect 193340 140588 193396 140644
rect 192780 140476 192836 140532
rect 191996 140364 192052 140420
rect 190988 140252 191044 140308
rect 185724 140140 185780 140196
rect 190988 139916 191044 139972
rect 191996 140028 192052 140084
rect 192780 139468 192836 139524
rect 193340 140252 193396 140308
rect 196700 139132 196756 139188
rect 185612 138796 185668 138852
rect 225148 153692 225204 153748
rect 230300 156492 230356 156548
rect 234332 156492 234388 156548
rect 232988 145740 233044 145796
rect 233100 147084 233156 147140
rect 227612 145628 227668 145684
rect 222572 143948 222628 144004
rect 224924 143948 224980 144004
rect 212940 142380 212996 142436
rect 223804 141484 223860 141540
rect 214620 141148 214676 141204
rect 219324 141148 219380 141204
rect 217420 140812 217476 140868
rect 216412 140476 216468 140532
rect 216412 139804 216468 139860
rect 217420 140364 217476 140420
rect 223356 139356 223412 139412
rect 234332 143948 234388 144004
rect 235676 143612 235732 143668
rect 235788 150444 235844 150500
rect 241948 157164 242004 157220
rect 246428 157164 246484 157220
rect 247772 157388 247828 157444
rect 246652 157052 246708 157108
rect 243740 156268 243796 156324
rect 246092 156268 246148 156324
rect 241948 150668 242004 150724
rect 241052 145516 241108 145572
rect 243852 146972 243908 147028
rect 238364 145404 238420 145460
rect 235004 142268 235060 142324
rect 234556 141820 234612 141876
rect 234220 141372 234276 141428
rect 233772 139580 233828 139636
rect 233996 139132 234052 139188
rect 235004 141820 235060 141876
rect 235116 142156 235172 142212
rect 235116 141372 235172 141428
rect 235004 139244 235060 139300
rect 249116 157052 249172 157108
rect 251804 156268 251860 156324
rect 252812 157500 252868 157556
rect 247772 147420 247828 147476
rect 249340 148652 249396 148708
rect 246652 147196 246708 147252
rect 246092 143724 246148 143780
rect 247548 146188 247604 146244
rect 244636 141148 244692 141204
rect 245420 140588 245476 140644
rect 223356 138908 223412 138964
rect 196924 138796 196980 138852
rect 218204 138684 218260 138740
rect 234780 138572 234836 138628
rect 195916 39452 195972 39508
rect 176988 14252 177044 14308
rect 160860 4620 160916 4676
rect 175084 4620 175140 4676
rect 163884 4508 163940 4564
rect 161980 4396 162036 4452
rect 169596 4284 169652 4340
rect 167916 4172 167972 4228
rect 165788 4060 165844 4116
rect 171388 4172 171444 4228
rect 173404 3836 173460 3892
rect 184604 12572 184660 12628
rect 182924 6076 182980 6132
rect 179116 4060 179172 4116
rect 181020 4060 181076 4116
rect 186732 7644 186788 7700
rect 190540 7532 190596 7588
rect 188636 4060 188692 4116
rect 192444 4284 192500 4340
rect 194348 4172 194404 4228
rect 197932 37884 197988 37940
rect 195916 4172 195972 4228
rect 196028 37772 196084 37828
rect 209356 36204 209412 36260
rect 201740 36092 201796 36148
rect 199948 29372 200004 29428
rect 207452 32732 207508 32788
rect 203644 31052 203700 31108
rect 205772 4396 205828 4452
rect 221004 5964 221060 6020
rect 215292 5852 215348 5908
rect 211484 4508 211540 4564
rect 238140 4620 238196 4676
rect 226716 4060 226772 4116
rect 232428 4060 232484 4116
rect 247548 4284 247604 4340
rect 243852 4172 243908 4228
rect 257180 159404 257236 159460
rect 260428 158844 260484 158900
rect 262556 157836 262612 157892
rect 265244 157500 265300 157556
rect 254492 157276 254548 157332
rect 265468 157276 265524 157332
rect 261212 157164 261268 157220
rect 258636 156268 258692 156324
rect 258636 155596 258692 155652
rect 252812 147084 252868 147140
rect 255052 152348 255108 152404
rect 250348 143836 250404 143892
rect 250348 4172 250404 4228
rect 257852 151116 257908 151172
rect 260316 148764 260372 148820
rect 257852 4508 257908 4564
rect 259532 138908 259588 138964
rect 259532 4396 259588 4452
rect 264572 157052 264628 157108
rect 270620 157724 270676 157780
rect 273868 158844 273924 158900
rect 273868 157836 273924 157892
rect 277676 158956 277732 159012
rect 275996 157836 276052 157892
rect 273308 157612 273364 157668
rect 267932 157052 267988 157108
rect 265468 150444 265524 150500
rect 279132 301420 279188 301476
rect 294812 352492 294868 352548
rect 293132 324268 293188 324324
rect 289772 266364 289828 266420
rect 291452 322924 291508 322980
rect 284732 170492 284788 170548
rect 293132 163772 293188 163828
rect 291452 162092 291508 162148
rect 279132 160300 279188 160356
rect 279020 160188 279076 160244
rect 278908 152348 278964 152404
rect 278796 148652 278852 148708
rect 284284 152236 284340 152292
rect 273420 147420 273476 147476
rect 264572 146972 264628 147028
rect 265356 147308 265412 147364
rect 261212 143836 261268 143892
rect 263788 141932 263844 141988
rect 264460 141820 264516 141876
rect 264460 141260 264516 141316
rect 276108 144060 276164 144116
rect 274988 141708 275044 141764
rect 274540 141596 274596 141652
rect 274204 139692 274260 139748
rect 274988 141372 275044 141428
rect 263788 138908 263844 138964
rect 275436 139020 275492 139076
rect 296492 372652 296548 372708
rect 388892 368732 388948 368788
rect 299852 353836 299908 353892
rect 296492 273084 296548 273140
rect 298172 329644 298228 329700
rect 294924 264796 294980 264852
rect 299852 271628 299908 271684
rect 298172 168812 298228 168868
rect 294812 152236 294868 152292
rect 285068 142044 285124 142100
rect 285068 141260 285124 141316
rect 308252 275660 308308 275716
rect 304444 269948 304500 270004
rect 308252 215964 308308 216020
rect 309932 275548 309988 275604
rect 313292 275548 313348 275604
rect 309932 214284 309988 214340
rect 308252 157052 308308 157108
rect 308252 156156 308308 156212
rect 306572 155708 306628 155764
rect 304780 142716 304836 142772
rect 303212 140588 303268 140644
rect 293356 140252 293412 140308
rect 285740 140140 285796 140196
rect 292012 140028 292068 140084
rect 285740 139804 285796 139860
rect 291004 139916 291060 139972
rect 292012 139580 292068 139636
rect 292796 140028 292852 140084
rect 292796 139468 292852 139524
rect 293356 139468 293412 139524
rect 312508 142940 312564 142996
rect 314076 142940 314132 142996
rect 315420 144060 315476 144116
rect 315420 143164 315476 143220
rect 312508 139244 312564 139300
rect 312956 142380 313012 142436
rect 314636 141148 314692 141204
rect 315532 143276 315588 143332
rect 315868 275660 315924 275716
rect 329644 275548 329700 275604
rect 322588 222684 322644 222740
rect 330876 276332 330932 276388
rect 330876 275548 330932 275604
rect 315756 144060 315812 144116
rect 315756 143052 315812 143108
rect 324940 155820 324996 155876
rect 315756 142268 315812 142324
rect 316428 142268 316484 142324
rect 315532 142156 315588 142212
rect 315420 139132 315476 139188
rect 316428 140476 316484 140532
rect 317436 142044 317492 142100
rect 317436 140364 317492 140420
rect 318220 141708 318276 141764
rect 319228 141148 319284 141204
rect 323596 139244 323652 139300
rect 323820 142380 323876 142436
rect 323820 141484 323876 141540
rect 325052 142380 325108 142436
rect 330316 262668 330372 262724
rect 332444 262892 332500 262948
rect 330876 142716 330932 142772
rect 331772 262108 331828 262164
rect 331772 142268 331828 142324
rect 330316 141708 330372 141764
rect 330876 141708 330932 141764
rect 332556 262108 332612 262164
rect 332444 142044 332500 142100
rect 333116 150556 333172 150612
rect 331772 140924 331828 140980
rect 330876 139132 330932 139188
rect 334124 143276 334180 143332
rect 333452 142716 333508 142772
rect 333788 143164 333844 143220
rect 296828 138796 296884 138852
rect 317772 138684 317828 138740
rect 334124 141932 334180 141988
rect 342636 215852 342692 215908
rect 347788 279804 347844 279860
rect 335692 150668 335748 150724
rect 334348 142828 334404 142884
rect 334348 141708 334404 141764
rect 334572 143052 334628 143108
rect 334572 141484 334628 141540
rect 335020 142940 335076 142996
rect 335020 140588 335076 140644
rect 343868 147196 343924 147252
rect 336028 142044 336084 142100
rect 336028 140140 336084 140196
rect 344652 142044 344708 142100
rect 345324 141148 345380 141204
rect 345324 139020 345380 139076
rect 333788 138684 333844 138740
rect 275324 138572 275380 138628
rect 260316 4172 260372 4228
rect 260764 14252 260820 14308
rect 317884 7532 317940 7588
rect 295036 5964 295092 6020
rect 283612 5068 283668 5124
rect 266700 4284 266756 4340
rect 272188 4172 272244 4228
rect 277900 4172 277956 4228
rect 289324 5068 289380 5124
rect 312172 5964 312228 6020
rect 300748 5068 300804 5124
rect 306460 4172 306516 4228
rect 346668 4284 346724 4340
rect 323596 4172 323652 4228
rect 329308 4172 329364 4228
rect 335244 4172 335300 4228
rect 340956 4172 341012 4228
rect 347900 278348 347956 278404
rect 350252 276780 350308 276836
rect 347900 4508 347956 4564
rect 348012 273196 348068 273252
rect 350252 212492 350308 212548
rect 350476 276556 350532 276612
rect 355292 279692 355348 279748
rect 352044 275548 352100 275604
rect 353948 275548 354004 275604
rect 353612 269836 353668 269892
rect 350476 4956 350532 5012
rect 352156 168812 352212 168868
rect 348012 4284 348068 4340
rect 347788 4172 347844 4228
rect 353948 269836 354004 269892
rect 353612 20300 353668 20356
rect 356748 268268 356804 268324
rect 356076 266588 356132 266644
rect 363804 275548 363860 275604
rect 363132 273196 363188 273252
rect 359436 269948 359492 270004
rect 364588 268156 364644 268212
rect 366268 275548 366324 275604
rect 366268 268156 366324 268212
rect 364476 266700 364532 266756
rect 357756 265020 357812 265076
rect 363804 265132 363860 265188
rect 357084 262780 357140 262836
rect 355292 4844 355348 4900
rect 356972 257852 357028 257908
rect 360332 262444 360388 262500
rect 364252 259084 364308 259140
rect 374108 278796 374164 278852
rect 374444 278796 374500 278852
rect 371308 266476 371364 266532
rect 365372 262780 365428 262836
rect 373772 262780 373828 262836
rect 373436 262444 373492 262500
rect 374556 263004 374612 263060
rect 374332 262444 374388 262500
rect 374556 262780 374612 262836
rect 374220 262220 374276 262276
rect 373884 258972 373940 259028
rect 375452 276780 375508 276836
rect 380492 275660 380548 275716
rect 380492 266700 380548 266756
rect 382172 275548 382228 275604
rect 384412 275660 384468 275716
rect 383516 275548 383572 275604
rect 383852 275548 383908 275604
rect 385196 275548 385252 275604
rect 385308 273196 385364 273252
rect 383852 265132 383908 265188
rect 385084 268156 385140 268212
rect 382172 264908 382228 264964
rect 375452 263004 375508 263060
rect 374668 262220 374724 262276
rect 375004 262444 375060 262500
rect 375004 259084 375060 259140
rect 376124 262108 376180 262164
rect 363916 258636 363972 258692
rect 374332 258636 374388 258692
rect 384300 258860 384356 258916
rect 419132 342748 419188 342804
rect 460236 418124 460292 418180
rect 460124 416556 460180 416612
rect 456092 276668 456148 276724
rect 459452 381388 459508 381444
rect 419356 276332 419412 276388
rect 388892 262556 388948 262612
rect 390572 269948 390628 270004
rect 385756 259084 385812 259140
rect 396844 269836 396900 269892
rect 392812 268268 392868 268324
rect 391916 265020 391972 265076
rect 390572 259084 390628 259140
rect 392252 258972 392308 259028
rect 393372 266588 393428 266644
rect 393932 259084 393988 259140
rect 417452 262892 417508 262948
rect 416332 262332 416388 262388
rect 397292 259084 397348 259140
rect 418124 262668 418180 262724
rect 454972 271628 455028 271684
rect 423948 261324 424004 261380
rect 435708 260428 435764 260484
rect 432236 259756 432292 259812
rect 443436 259644 443492 259700
rect 392476 258972 392532 259028
rect 385420 258860 385476 258916
rect 406588 258748 406644 258804
rect 412412 258748 412468 258804
rect 414092 258748 414148 258804
rect 424396 258748 424452 258804
rect 375228 258636 375284 258692
rect 434924 258636 434980 258692
rect 433804 258524 433860 258580
rect 423388 258412 423444 258468
rect 434140 258412 434196 258468
rect 434588 258412 434644 258468
rect 444668 258412 444724 258468
rect 445340 258412 445396 258468
rect 360332 254492 360388 254548
rect 357084 217644 357140 217700
rect 356972 4060 357028 4116
rect 357868 170492 357924 170548
rect 443884 155484 443940 155540
rect 406588 155372 406644 155428
rect 384412 153692 384468 153748
rect 365372 145740 365428 145796
rect 364252 142268 364308 142324
rect 364476 142268 364532 142324
rect 364476 141820 364532 141876
rect 376124 145628 376180 145684
rect 373436 143948 373492 144004
rect 373324 141820 373380 141876
rect 373324 141372 373380 141428
rect 374556 142156 374612 142212
rect 374556 141148 374612 141204
rect 374220 139692 374276 139748
rect 375004 141820 375060 141876
rect 375452 141372 375508 141428
rect 385084 141260 385140 141316
rect 391916 140812 391972 140868
rect 391020 140252 391076 140308
rect 391020 139916 391076 139972
rect 385756 139804 385812 139860
rect 393372 140700 393428 140756
rect 391916 139580 391972 139636
rect 392812 140476 392868 140532
rect 392812 140028 392868 140084
rect 393372 139468 393428 139524
rect 424956 152124 425012 152180
rect 412412 142716 412468 142772
rect 412412 141708 412468 141764
rect 423724 142380 423780 142436
rect 423724 141820 423780 141876
rect 414652 141148 414708 141204
rect 419244 141148 419300 141204
rect 416332 140924 416388 140980
rect 417452 140140 417508 140196
rect 417676 139132 417732 139188
rect 423612 139132 423668 139188
rect 433132 150332 433188 150388
rect 435708 147084 435764 147140
rect 434140 141932 434196 141988
rect 433804 141708 433860 141764
rect 433804 140028 433860 140084
rect 363804 138908 363860 138964
rect 418124 138908 418180 138964
rect 396844 138796 396900 138852
rect 434588 141484 434644 141540
rect 434812 140588 434868 140644
rect 433804 138684 433860 138740
rect 449260 152236 449316 152292
rect 444668 141932 444724 141988
rect 445564 139020 445620 139076
rect 434924 138684 434980 138740
rect 375228 138572 375284 138628
rect 437836 36092 437892 36148
rect 426412 17612 426468 17668
rect 420700 15932 420756 15988
rect 392140 14252 392196 14308
rect 363580 4956 363636 5012
rect 375004 4844 375060 4900
rect 369292 4060 369348 4116
rect 380716 4732 380772 4788
rect 386428 4620 386484 4676
rect 409276 5852 409332 5908
rect 403564 4508 403620 4564
rect 397852 4396 397908 4452
rect 414988 4284 415044 4340
rect 432124 4172 432180 4228
rect 443772 4172 443828 4228
rect 460124 37772 460180 37828
rect 462812 432796 462868 432852
rect 462924 555212 462980 555268
rect 461244 432684 461300 432740
rect 461132 377804 461188 377860
rect 462812 430108 462868 430164
rect 474348 583772 474404 583828
rect 518476 590940 518532 590996
rect 496412 582204 496468 582260
rect 540540 582092 540596 582148
rect 584668 591276 584724 591332
rect 562604 578732 562660 578788
rect 464492 444444 464548 444500
rect 464604 555324 464660 555380
rect 468524 551516 468580 551572
rect 468412 551404 468468 551460
rect 468300 551292 468356 551348
rect 468188 551180 468244 551236
rect 467740 549500 467796 549556
rect 468076 549052 468132 549108
rect 467740 501564 467796 501620
rect 467852 548268 467908 548324
rect 467740 495516 467796 495572
rect 467964 546924 468020 546980
rect 468076 465276 468132 465332
rect 468188 507612 468244 507668
rect 467964 459228 468020 459284
rect 467852 453180 467908 453236
rect 467740 450380 467796 450436
rect 464604 432908 464660 432964
rect 468300 513660 468356 513716
rect 468412 519708 468468 519764
rect 468524 525756 468580 525812
rect 468636 549388 468692 549444
rect 495516 537740 495572 537796
rect 468636 531804 468692 531860
rect 470316 537628 470372 537684
rect 470092 500892 470148 500948
rect 468636 446796 468692 446852
rect 469868 459228 469924 459284
rect 468524 397740 468580 397796
rect 468636 421260 468692 421316
rect 468412 396172 468468 396228
rect 468300 394604 468356 394660
rect 468188 393036 468244 393092
rect 462924 377692 462980 377748
rect 467852 377132 467908 377188
rect 467852 160636 467908 160692
rect 469980 403340 470036 403396
rect 470092 391468 470148 391524
rect 470204 464604 470260 464660
rect 469980 386764 470036 386820
rect 477596 537628 477652 537684
rect 547148 537628 547204 537684
rect 512316 535948 512372 536004
rect 554428 537628 554484 537684
rect 529340 534268 529396 534324
rect 470316 451500 470372 451556
rect 470652 452396 470708 452452
rect 470204 385196 470260 385252
rect 469868 383628 469924 383684
rect 474908 450492 474964 450548
rect 470876 450380 470932 450436
rect 470876 389900 470932 389956
rect 472892 450268 472948 450324
rect 533036 450156 533092 450212
rect 474908 448364 474964 448420
rect 479612 448364 479668 448420
rect 477932 447916 477988 447972
rect 475132 447692 475188 447748
rect 474572 446796 474628 446852
rect 474572 399308 474628 399364
rect 477596 429772 477652 429828
rect 477036 422828 477092 422884
rect 476924 419692 476980 419748
rect 476252 414988 476308 415044
rect 476252 402892 476308 402948
rect 476476 413420 476532 413476
rect 476476 402780 476532 402836
rect 475132 398076 475188 398132
rect 472892 388332 472948 388388
rect 476252 397292 476308 397348
rect 470652 382060 470708 382116
rect 476252 334796 476308 334852
rect 476364 383852 476420 383908
rect 476924 379036 476980 379092
rect 477596 402220 477652 402276
rect 477820 429660 477876 429716
rect 478492 447804 478548 447860
rect 478044 443212 478100 443268
rect 478380 432012 478436 432068
rect 478044 402332 478100 402388
rect 478156 431900 478212 431956
rect 477932 401436 477988 401492
rect 478380 402556 478436 402612
rect 478156 401324 478212 401380
rect 478716 425964 478772 426020
rect 478492 399756 478548 399812
rect 478604 424396 478660 424452
rect 477820 399644 477876 399700
rect 477036 375452 477092 375508
rect 477932 377356 477988 377412
rect 476364 333900 476420 333956
rect 476476 325836 476532 325892
rect 476252 324940 476308 324996
rect 476140 312396 476196 312452
rect 476140 293916 476196 293972
rect 476364 322252 476420 322308
rect 476700 324044 476756 324100
rect 476476 300524 476532 300580
rect 476588 314188 476644 314244
rect 476364 297164 476420 297220
rect 476252 292236 476308 292292
rect 476924 323148 476980 323204
rect 476700 300636 476756 300692
rect 476812 316876 476868 316932
rect 476924 302316 476980 302372
rect 477036 315980 477092 316036
rect 476812 297276 476868 297332
rect 476588 290556 476644 290612
rect 477036 288988 477092 289044
rect 478604 373772 478660 373828
rect 480620 446908 480676 446964
rect 479612 379372 479668 379428
rect 480060 426860 480116 426916
rect 478716 372092 478772 372148
rect 479612 377244 479668 377300
rect 484092 446908 484148 446964
rect 488124 449596 488180 449652
rect 482748 444444 482804 444500
rect 485436 432908 485492 432964
rect 484092 432796 484148 432852
rect 486780 432684 486836 432740
rect 493500 447916 493556 447972
rect 502908 447804 502964 447860
rect 504252 449484 504308 449540
rect 489468 437836 489524 437892
rect 490812 432572 490868 432628
rect 497532 432236 497588 432292
rect 496188 432124 496244 432180
rect 492156 432012 492212 432068
rect 494844 431900 494900 431956
rect 493500 431788 493556 431844
rect 498876 432124 498932 432180
rect 502908 432012 502964 432068
rect 512316 447692 512372 447748
rect 521612 448476 521668 448532
rect 527436 449372 527492 449428
rect 527436 448476 527492 448532
rect 531132 448476 531188 448532
rect 521612 447356 521668 447412
rect 525756 447804 525812 447860
rect 509628 446124 509684 446180
rect 506940 444332 506996 444388
rect 505596 434364 505652 434420
rect 508284 437724 508340 437780
rect 510972 434252 511028 434308
rect 512316 432572 512372 432628
rect 519036 431900 519092 431956
rect 513660 429884 513716 429940
rect 523068 431788 523124 431844
rect 521724 430220 521780 430276
rect 519596 429996 519652 430052
rect 524412 430108 524468 430164
rect 527100 447692 527156 447748
rect 532700 446012 532756 446068
rect 532588 439292 532644 439348
rect 515004 429772 515060 429828
rect 516348 429660 516404 429716
rect 517692 429436 517748 429492
rect 500220 429324 500276 429380
rect 501564 429212 501620 429268
rect 532588 426412 532644 426468
rect 532700 421036 532756 421092
rect 532812 437612 532868 437668
rect 532812 415660 532868 415716
rect 532924 429548 532980 429604
rect 532924 410284 532980 410340
rect 480620 400204 480676 400260
rect 540540 447804 540596 447860
rect 549948 447692 550004 447748
rect 533372 407372 533428 407428
rect 557788 508284 557844 508340
rect 557788 451276 557844 451332
rect 557900 497756 557956 497812
rect 557900 451164 557956 451220
rect 558012 487228 558068 487284
rect 590492 482860 590548 482916
rect 558124 476700 558180 476756
rect 558124 451388 558180 451444
rect 558236 466172 558292 466228
rect 558236 451052 558292 451108
rect 590492 450492 590548 450548
rect 558012 450268 558068 450324
rect 554428 407372 554484 407428
rect 533372 404908 533428 404964
rect 533372 390572 533428 390628
rect 533372 388780 533428 388836
rect 533036 383404 533092 383460
rect 484764 380716 484820 380772
rect 590604 380492 590660 380548
rect 502908 380380 502964 380436
rect 526316 380380 526372 380436
rect 500892 380268 500948 380324
rect 482748 380156 482804 380212
rect 488796 377804 488852 377860
rect 486780 377692 486836 377748
rect 492828 380044 492884 380100
rect 496860 379484 496916 379540
rect 494844 377916 494900 377972
rect 498876 377916 498932 377972
rect 490812 377580 490868 377636
rect 504924 377468 504980 377524
rect 480060 368844 480116 368900
rect 508956 377356 509012 377412
rect 510972 377244 511028 377300
rect 515004 379372 515060 379428
rect 519036 379596 519092 379652
rect 517020 378924 517076 378980
rect 523068 380044 523124 380100
rect 521052 377916 521108 377972
rect 525084 377916 525140 377972
rect 559468 379036 559524 379092
rect 512988 377132 513044 377188
rect 506940 368732 506996 368788
rect 482524 348572 482580 348628
rect 498988 345324 499044 345380
rect 495964 344876 496020 344932
rect 492604 344652 492660 344708
rect 482524 342748 482580 342804
rect 485884 344540 485940 344596
rect 489244 344428 489300 344484
rect 502348 345324 502404 345380
rect 505708 345324 505764 345380
rect 509404 344428 509460 344484
rect 512764 344428 512820 344484
rect 516124 344428 516180 344484
rect 519484 344428 519540 344484
rect 479612 271516 479668 271572
rect 477932 266252 477988 266308
rect 468636 158956 468692 159012
rect 464716 155372 464772 155428
rect 462812 149660 462868 149716
rect 464492 150332 464548 150388
rect 463820 142716 463876 142772
rect 463820 142044 463876 142100
rect 464716 142716 464772 142772
rect 465388 150444 465444 150500
rect 464492 142268 464548 142324
rect 475020 159404 475076 159460
rect 483980 159628 484036 159684
rect 483196 158732 483252 158788
rect 474572 156268 474628 156324
rect 472892 141932 472948 141988
rect 473452 155596 473508 155652
rect 474572 152124 474628 152180
rect 474124 147084 474180 147140
rect 474124 141148 474180 141204
rect 475468 150444 475524 150500
rect 474572 142156 474628 142212
rect 475020 145628 475076 145684
rect 475020 142492 475076 142548
rect 476028 146972 476084 147028
rect 484092 141708 484148 141764
rect 484316 143836 484372 143892
rect 485212 159628 485268 159684
rect 484652 142044 484708 142100
rect 485100 143836 485156 143892
rect 485100 142604 485156 142660
rect 484764 140588 484820 140644
rect 484764 140028 484820 140084
rect 484876 141708 484932 141764
rect 485884 158844 485940 158900
rect 493948 157500 494004 157556
rect 501228 160076 501284 160132
rect 493052 155596 493108 155652
rect 491372 155484 491428 155540
rect 485436 141708 485492 141764
rect 486332 152236 486388 152292
rect 486332 140364 486388 140420
rect 491372 140252 491428 140308
rect 491596 150556 491652 150612
rect 491596 140812 491652 140868
rect 493052 140476 493108 140532
rect 493388 146972 493444 147028
rect 494732 141820 494788 141876
rect 495404 142940 495460 142996
rect 493388 140700 493444 140756
rect 496860 145740 496916 145796
rect 495516 142156 495572 142212
rect 495516 141820 495572 141876
rect 495404 139132 495460 139188
rect 500556 142828 500612 142884
rect 498988 142268 499044 142324
rect 502124 160076 502180 160132
rect 501452 142268 501508 142324
rect 498988 140140 499044 140196
rect 500668 141260 500724 141316
rect 502236 141260 502292 141316
rect 505596 141484 505652 141540
rect 506604 152012 506660 152068
rect 503916 141372 503972 141428
rect 503916 140924 503972 140980
rect 500668 139132 500724 139188
rect 496860 139020 496916 139076
rect 512316 159516 512372 159572
rect 526092 155596 526148 155652
rect 527996 155484 528052 155540
rect 533148 152236 533204 152292
rect 526988 150556 527044 150612
rect 542892 157724 542948 157780
rect 534604 156156 534660 156212
rect 542556 150444 542612 150500
rect 544348 152124 544404 152180
rect 524188 146972 524244 147028
rect 520828 145740 520884 145796
rect 545468 157612 545524 157668
rect 552076 158956 552132 159012
rect 544572 147084 544628 147140
rect 542668 145628 542724 145684
rect 532588 143836 532644 143892
rect 533036 145516 533092 145572
rect 524972 143724 525028 143780
rect 523404 142940 523460 142996
rect 519260 142828 519316 142884
rect 517468 142268 517524 142324
rect 507276 141596 507332 141652
rect 512988 141596 513044 141652
rect 514668 141484 514724 141540
rect 516348 141372 516404 141428
rect 518140 141260 518196 141316
rect 523740 142156 523796 142212
rect 535724 145404 535780 145460
rect 534156 142044 534212 142100
rect 533820 140588 533876 140644
rect 534940 141708 534996 141764
rect 534604 141148 534660 141204
rect 543900 143612 543956 143668
rect 545356 141932 545412 141988
rect 544684 141148 544740 141204
rect 484876 138684 484932 138740
rect 475244 138572 475300 138628
rect 460236 36092 460292 36148
rect 460684 39452 460740 39508
rect 459452 4172 459508 4228
rect 489244 37996 489300 38052
rect 466396 5964 466452 6020
rect 472108 4620 472164 4676
rect 477820 4508 477876 4564
rect 483532 4396 483588 4452
rect 512092 37884 512148 37940
rect 506380 24332 506436 24388
rect 500668 5852 500724 5908
rect 494956 4284 495012 4340
rect 534940 37772 534996 37828
rect 517804 34412 517860 34468
rect 529228 32732 529284 32788
rect 523516 4172 523572 4228
rect 540652 36092 540708 36148
rect 546588 4172 546644 4228
rect 553532 157836 553588 157892
rect 555100 155372 555156 155428
rect 554316 150332 554372 150388
rect 590492 378812 590548 378868
rect 559468 4284 559524 4340
rect 559580 375452 559636 375508
rect 558012 4172 558068 4228
rect 559580 4172 559636 4228
rect 563500 373772 563556 373828
rect 569212 372092 569268 372148
rect 565292 278236 565348 278292
rect 568652 269612 568708 269668
rect 568652 139244 568708 139300
rect 565292 7084 565348 7140
rect 574924 368844 574980 368900
rect 570332 276444 570388 276500
rect 570332 178892 570388 178948
rect 590604 364140 590660 364196
rect 590492 324492 590548 324548
rect 590604 278124 590660 278180
rect 580636 273084 580692 273140
rect 582540 266364 582596 266420
rect 584444 264796 584500 264852
rect 590492 264572 590548 264628
rect 590716 268044 590772 268100
rect 590716 245196 590772 245252
rect 590604 165900 590660 165956
rect 590604 160412 590660 160468
rect 590604 86604 590660 86660
rect 590492 46956 590548 47012
<< metal3 >>
rect 320114 591276 320124 591332
rect 320180 591276 464492 591332
rect 464548 591276 464558 591332
rect 584658 591276 584668 591332
rect 584724 591276 584762 591332
rect 298050 591164 298060 591220
rect 298116 591164 451276 591220
rect 451332 591164 451342 591220
rect 231746 591052 231756 591108
rect 231812 591052 449372 591108
rect 449428 591052 449438 591108
rect 209794 590940 209804 590996
rect 209860 590940 279692 590996
rect 279748 590940 279758 590996
rect 299954 590940 299964 590996
rect 300020 590940 518476 590996
rect 518532 590940 518542 590996
rect 165666 590828 165676 590884
rect 165732 590828 456204 590884
rect 456260 590828 456270 590884
rect 99474 590716 99484 590772
rect 99540 590716 457772 590772
rect 457828 590716 457838 590772
rect 55346 590604 55356 590660
rect 55412 590604 459564 590660
rect 459620 590604 459630 590660
rect 33282 590492 33292 590548
rect 33348 590492 451052 590548
rect 451108 590492 451118 590548
rect 298274 590380 298284 590436
rect 298340 590380 386092 590436
rect 386148 590380 386158 590436
rect 275986 590156 275996 590212
rect 276052 590156 278012 590212
rect 278068 590156 278078 590212
rect 253922 588924 253932 588980
rect 253988 588924 462812 588980
rect 462868 588924 462878 588980
rect 50306 588812 50316 588868
rect 50372 588812 408268 588868
rect 408324 588812 408334 588868
rect 595560 588644 597000 588840
rect 51986 588588 51996 588644
rect 52052 588616 597000 588644
rect 52052 588588 595672 588616
rect -960 587188 480 587384
rect -960 587160 456092 587188
rect 392 587132 456092 587160
rect 456148 587132 456158 587188
rect 55346 583772 55356 583828
rect 55412 583772 474348 583828
rect 474404 583772 474414 583828
rect 58706 582204 58716 582260
rect 58772 582204 496412 582260
rect 496468 582204 496478 582260
rect 53666 582092 53676 582148
rect 53732 582092 540540 582148
rect 540596 582092 540606 582148
rect 51874 578732 51884 578788
rect 51940 578732 562604 578788
rect 562660 578732 562670 578788
rect 595560 575428 597000 575624
rect 50306 575372 50316 575428
rect 50372 575400 597000 575428
rect 50372 575372 595672 575400
rect -960 573076 480 573272
rect -960 573048 452732 573076
rect 392 573020 452732 573048
rect 452788 573020 452798 573076
rect 58482 572124 58492 572180
rect 58548 572124 341964 572180
rect 342020 572124 342030 572180
rect 121762 572012 121772 572068
rect 121828 572012 452284 572068
rect 452340 572012 452350 572068
rect 121314 570332 121324 570388
rect 121380 570332 461244 570388
rect 461300 570332 461310 570388
rect 57026 566972 57036 567028
rect 57092 566972 364028 567028
rect 364084 566972 364094 567028
rect 58594 565404 58604 565460
rect 58660 565404 430220 565460
rect 430276 565404 430286 565460
rect 77298 565292 77308 565348
rect 77364 565292 461132 565348
rect 461188 565292 461198 565348
rect 10994 563612 11004 563668
rect 11060 563612 454412 563668
rect 454468 563612 454478 563668
rect 595560 562212 597000 562408
rect 279794 562156 279804 562212
rect 279860 562184 597000 562212
rect 279860 562156 595672 562184
rect -960 558964 480 559160
rect -960 558936 4172 558964
rect 392 558908 4172 558936
rect 4228 558908 4238 558964
rect 153682 557788 153692 557844
rect 153748 557788 173740 557844
rect 173796 557788 173806 557844
rect 187506 555324 187516 555380
rect 187572 555324 464604 555380
rect 464660 555324 464670 555380
rect 143378 555212 143388 555268
rect 143444 555212 462924 555268
rect 462980 555212 462990 555268
rect 274642 554428 274652 554484
rect 274708 554428 416780 554484
rect 416836 554428 416846 554484
rect 201282 554316 201292 554372
rect 201348 554316 212492 554372
rect 212548 554316 212558 554372
rect 278114 553532 278124 553588
rect 278180 553532 426636 553588
rect 426692 553532 426702 553588
rect 291442 553420 291452 553476
rect 291508 553420 421708 553476
rect 421764 553420 421774 553476
rect 318210 553308 318220 553364
rect 318276 553308 452844 553364
rect 452900 553308 452910 553364
rect 313282 553196 313292 553252
rect 313348 553196 451164 553252
rect 451220 553196 451230 553252
rect 303426 553084 303436 553140
rect 303492 553084 449484 553140
rect 449540 553084 449550 553140
rect 308354 552972 308364 553028
rect 308420 552972 454524 553028
rect 454580 552972 454590 553028
rect 289762 552860 289772 552916
rect 289828 552860 436492 552916
rect 436548 552860 436558 552916
rect 214872 551516 216748 551572
rect 216804 551516 216814 551572
rect 382386 551516 382396 551572
rect 382452 551516 468524 551572
rect 468580 551516 468590 551572
rect 377346 551404 377356 551460
rect 377412 551404 468412 551460
rect 468468 551404 468478 551460
rect 372418 551292 372428 551348
rect 372484 551292 468300 551348
rect 468356 551292 468366 551348
rect 367490 551180 367500 551236
rect 367556 551180 468188 551236
rect 468244 551180 468254 551236
rect 299842 551068 299852 551124
rect 299908 551068 406924 551124
rect 406980 551068 406990 551124
rect 217522 550172 217532 550228
rect 217588 550172 377356 550228
rect 377412 550172 377422 550228
rect 301074 550060 301084 550116
rect 301140 550060 430780 550116
rect 430836 550060 430846 550116
rect 301746 549948 301756 550004
rect 301812 549948 367164 550004
rect 367220 549948 367230 550004
rect 301858 549836 301868 549892
rect 301924 549836 372428 549892
rect 372484 549836 372494 549892
rect 384692 549836 397068 549892
rect 397124 549836 397134 549892
rect 384692 549780 384748 549836
rect 296482 549724 296492 549780
rect 296548 549724 384748 549780
rect 387174 549724 387212 549780
rect 387268 549724 392812 549780
rect 392868 549724 392878 549780
rect 293122 549612 293132 549668
rect 293188 549612 411852 549668
rect 411908 549612 411918 549668
rect 314132 549500 361228 549556
rect 362534 549500 362572 549556
rect 362628 549500 467740 549556
rect 467796 549500 467806 549556
rect 314132 549444 314188 549500
rect 361172 549444 361228 549500
rect 217746 549388 217756 549444
rect 217812 549388 314188 549444
rect 323110 549388 323148 549444
rect 323204 549388 323214 549444
rect 328038 549388 328076 549444
rect 328132 549388 328142 549444
rect 332966 549388 333004 549444
rect 333060 549388 333070 549444
rect 337894 549388 337932 549444
rect 337988 549388 337998 549444
rect 342822 549388 342860 549444
rect 342916 549388 342926 549444
rect 347750 549388 347788 549444
rect 347844 549388 347854 549444
rect 352678 549388 352716 549444
rect 352772 549388 352782 549444
rect 357606 549388 357644 549444
rect 357700 549388 357710 549444
rect 361172 549388 382284 549444
rect 382340 549388 382350 549444
rect 392102 549388 392140 549444
rect 392196 549388 392206 549444
rect 392802 549388 392812 549444
rect 392868 549388 468636 549444
rect 468692 549388 468702 549444
rect 294802 549276 294812 549332
rect 294868 549276 401996 549332
rect 402052 549276 402062 549332
rect 431330 549276 431340 549332
rect 431396 549276 431732 549332
rect 441410 549276 441420 549332
rect 441476 549276 459452 549332
rect 459508 549276 459518 549332
rect 431676 549220 431732 549276
rect 386978 549164 386988 549220
rect 387044 549164 392140 549220
rect 392196 549164 392206 549220
rect 431666 549164 431676 549220
rect 431732 549164 431742 549220
rect 301074 549052 301084 549108
rect 301140 549052 333004 549108
rect 333060 549052 468076 549108
rect 468132 549052 468142 549108
rect 595560 548996 597000 549192
rect 303426 548940 303436 548996
rect 303492 548940 342860 548996
rect 342916 548940 468300 548996
rect 468356 548940 468366 548996
rect 590146 548940 590156 548996
rect 590212 548968 597000 548996
rect 590212 548940 595672 548968
rect 214872 548828 215740 548884
rect 215796 548828 215806 548884
rect 300850 548828 300860 548884
rect 300916 548828 352716 548884
rect 352772 548828 468524 548884
rect 468580 548828 468590 548884
rect 298162 548716 298172 548772
rect 298228 548716 386988 548772
rect 387044 548716 387054 548772
rect 387202 548716 387212 548772
rect 387268 548716 387278 548772
rect 431666 548716 431676 548772
rect 431732 548716 446012 548772
rect 446068 548716 446078 548772
rect 387212 548660 387268 548716
rect 300962 548604 300972 548660
rect 301028 548604 387268 548660
rect 301634 548492 301644 548548
rect 301700 548492 362572 548548
rect 362628 548492 362638 548548
rect 303202 548380 303212 548436
rect 303268 548380 337932 548436
rect 337988 548380 337998 548436
rect 357634 548380 357644 548436
rect 357700 548380 467628 548436
rect 467684 548380 467694 548436
rect 323138 548268 323148 548324
rect 323204 548268 467852 548324
rect 467908 548268 467918 548324
rect 300962 547148 300972 547204
rect 301028 547148 323148 547204
rect 323204 547148 323214 547204
rect 301522 547036 301532 547092
rect 301588 547036 357644 547092
rect 357700 547036 357710 547092
rect 300738 546924 300748 546980
rect 300804 546924 328076 546980
rect 328132 546924 467964 546980
rect 468020 546924 468030 546980
rect 303314 546812 303324 546868
rect 303380 546812 347788 546868
rect 347844 546812 468188 546868
rect 468244 546812 468254 546868
rect 214872 546140 218428 546196
rect 218484 546140 218494 546196
rect 392 545048 4284 545076
rect -960 545020 4284 545048
rect 4340 545020 4350 545076
rect -960 544824 480 545020
rect 214872 543452 215180 543508
rect 215236 543452 215246 543508
rect 214872 540764 215292 540820
rect 215348 540764 215358 540820
rect 214872 538076 215404 538132
rect 215460 538076 215470 538132
rect 495506 537740 495516 537796
rect 495572 537740 548156 537796
rect 548212 537740 548222 537796
rect 470306 537628 470316 537684
rect 470372 537628 477596 537684
rect 477652 537628 477662 537684
rect 547138 537628 547148 537684
rect 547204 537628 554428 537684
rect 554484 537628 554494 537684
rect 512306 535948 512316 536004
rect 512372 535948 549388 536004
rect 549444 535948 549454 536004
rect 595560 535892 597000 535976
rect 590594 535836 590604 535892
rect 590660 535836 597000 535892
rect 595560 535752 597000 535836
rect 214872 535388 218540 535444
rect 218596 535388 218606 535444
rect 529302 534268 529340 534324
rect 529396 534268 529406 534324
rect 529330 533372 529340 533428
rect 529396 533372 549500 533428
rect 549556 533372 549566 533428
rect 214872 532700 217308 532756
rect 217364 532700 217374 532756
rect 468626 531804 468636 531860
rect 468692 531804 470120 531860
rect -960 530852 480 530936
rect -960 530796 4172 530852
rect 4228 530796 4238 530852
rect -960 530712 480 530796
rect 214872 530012 217084 530068
rect 217140 530012 300972 530068
rect 301028 530012 301038 530068
rect 554904 529340 556220 529396
rect 556276 529340 556286 529396
rect 214844 527436 217196 527492
rect 217252 527436 217756 527492
rect 217812 527436 217822 527492
rect 214844 527352 214900 527436
rect 468514 525756 468524 525812
rect 468580 525756 470120 525812
rect 214872 524636 217532 524692
rect 217588 524636 217598 524692
rect 590482 522732 590492 522788
rect 590548 522760 595672 522788
rect 590548 522732 597000 522760
rect 595560 522536 597000 522732
rect 214844 521668 214900 521976
rect 290612 521724 300524 521780
rect 300580 521724 300590 521780
rect 290612 521668 290668 521724
rect 214844 521612 216860 521668
rect 216916 521612 290668 521668
rect 297332 520268 300636 520324
rect 300692 520268 300702 520324
rect 297332 519988 297388 520268
rect 214844 519932 216972 519988
rect 217028 519932 297388 519988
rect 214844 519288 214900 519932
rect 468402 519708 468412 519764
rect 468468 519708 470120 519764
rect 554904 518812 556108 518868
rect 556164 518812 556174 518868
rect -960 516628 480 516824
rect 290612 516796 300524 516852
rect 300580 516796 300590 516852
rect 290612 516628 290668 516796
rect -960 516600 4284 516628
rect 392 516572 4284 516600
rect 4340 516572 4350 516628
rect 214872 516572 215516 516628
rect 215572 516572 290668 516628
rect 214872 513884 215628 513940
rect 215684 513884 215694 513940
rect 468290 513660 468300 513716
rect 468356 513660 470120 513716
rect 297332 513548 300636 513604
rect 300692 513548 300702 513604
rect 297332 513492 297388 513548
rect 290612 513436 297388 513492
rect 290612 513268 290668 513436
rect 215618 513212 215628 513268
rect 215684 513212 290668 513268
rect 214536 511224 300860 511252
rect 214508 511196 300860 511224
rect 300916 511196 300926 511252
rect 214508 510804 214564 511196
rect 214498 510748 214508 510804
rect 214564 510748 214574 510804
rect 595560 509348 597000 509544
rect 590706 509292 590716 509348
rect 590772 509320 597000 509348
rect 590772 509292 595672 509320
rect 214872 508536 215068 508564
rect 214844 508508 215068 508536
rect 215124 508508 215134 508564
rect 214844 508228 214900 508508
rect 554904 508284 557788 508340
rect 557844 508284 557854 508340
rect 214844 508172 301084 508228
rect 301140 508172 301150 508228
rect 468178 507612 468188 507668
rect 468244 507612 470120 507668
rect 214424 505848 300748 505876
rect 214396 505820 300748 505848
rect 300804 505820 300814 505876
rect 214396 505764 214452 505820
rect 214386 505708 214396 505764
rect 214452 505708 214462 505764
rect 214872 503160 300972 503188
rect 214844 503132 300972 503160
rect 301028 503132 301038 503188
rect 214844 502852 214900 503132
rect 214834 502796 214844 502852
rect 214900 502796 214910 502852
rect -960 502516 480 502712
rect -960 502488 4172 502516
rect 392 502460 4172 502488
rect 4228 502460 4238 502516
rect 176978 501676 176988 501732
rect 177044 501676 215404 501732
rect 215460 501676 215470 501732
rect 171490 501564 171500 501620
rect 171556 501564 217308 501620
rect 217364 501564 217374 501620
rect 467730 501564 467740 501620
rect 467796 501592 470120 501620
rect 467796 501564 470148 501592
rect 160850 501452 160860 501508
rect 160916 501452 215068 501508
rect 215124 501452 215134 501508
rect 470092 500948 470148 501564
rect 470082 500892 470092 500948
rect 470148 500892 470158 500948
rect 144722 500668 144732 500724
rect 144788 500668 217532 500724
rect 217588 500668 217598 500724
rect 176950 500556 176988 500612
rect 177044 500556 177054 500612
rect 171462 499996 171500 500052
rect 171556 499996 171566 500052
rect 155474 499884 155484 499940
rect 155540 499884 214844 499940
rect 214900 499884 214910 499940
rect 136658 499772 136668 499828
rect 136724 499772 215516 499828
rect 215572 499772 215582 499828
rect 150098 498204 150108 498260
rect 150164 498204 217084 498260
rect 217140 498204 217150 498260
rect 133970 498092 133980 498148
rect 134036 498092 215628 498148
rect 215684 498092 215694 498148
rect 554904 497756 557900 497812
rect 557956 497756 557966 497812
rect 202402 497196 202412 497252
rect 202468 497196 301084 497252
rect 301140 497196 301150 497252
rect 198594 496524 198604 496580
rect 198660 496524 284732 496580
rect 284788 496524 284798 496580
rect 194114 496412 194124 496468
rect 194180 496412 288092 496468
rect 288148 496412 288158 496468
rect 595560 496132 597000 496328
rect 590482 496076 590492 496132
rect 590548 496104 597000 496132
rect 590548 496076 595672 496104
rect 467618 495516 467628 495572
rect 467684 495516 467740 495572
rect 467796 495516 470120 495572
rect 147410 494732 147420 494788
rect 147476 494732 217196 494788
rect 217252 494732 217262 494788
rect 179666 493052 179676 493108
rect 179732 493052 215292 493108
rect 215348 493052 215358 493108
rect 182354 491372 182364 491428
rect 182420 491372 215180 491428
rect 215236 491372 215246 491428
rect 468626 489468 468636 489524
rect 468692 489468 470120 489524
rect -960 488404 480 488600
rect -960 488376 298396 488404
rect 392 488348 298396 488376
rect 298452 488348 298462 488404
rect 104402 488012 104412 488068
rect 104468 488012 299964 488068
rect 300020 488012 300030 488068
rect 554904 487228 558012 487284
rect 558068 487228 558078 487284
rect 20962 486332 20972 486388
rect 21028 486332 162764 486388
rect 162820 486332 162830 486388
rect 109778 484652 109788 484708
rect 109844 484652 298284 484708
rect 298340 484652 298350 484708
rect 468178 483420 468188 483476
rect 468244 483420 470120 483476
rect 595560 482916 597000 483112
rect 590482 482860 590492 482916
rect 590548 482888 597000 482916
rect 590548 482860 595672 482888
rect 468290 477372 468300 477428
rect 468356 477372 470120 477428
rect 554904 476700 558124 476756
rect 558180 476700 558190 476756
rect 63746 476252 63756 476308
rect 63812 476252 153692 476308
rect 153748 476252 153758 476308
rect -960 474292 480 474488
rect -960 474264 294924 474292
rect 392 474236 294924 474264
rect 294980 474236 294990 474292
rect 467842 471324 467852 471380
rect 467908 471324 470120 471380
rect 595560 469700 597000 469896
rect 590818 469644 590828 469700
rect 590884 469672 597000 469700
rect 590884 469644 595672 469672
rect 120530 469532 120540 469588
rect 120596 469532 212044 469588
rect 212100 469532 212110 469588
rect 22642 467852 22652 467908
rect 22708 467852 176204 467908
rect 176260 467852 176270 467908
rect 15922 466172 15932 466228
rect 15988 466172 189644 466228
rect 189700 466172 189710 466228
rect 554904 466172 558236 466228
rect 558292 466172 558302 466228
rect 468066 465276 468076 465332
rect 468132 465304 470232 465332
rect 468132 465276 470260 465304
rect 470204 464660 470260 465276
rect 470194 464604 470204 464660
rect 470260 464604 470270 464660
rect 14242 464492 14252 464548
rect 14308 464492 185164 464548
rect 185220 464492 185230 464548
rect -960 460180 480 460376
rect -960 460152 4396 460180
rect 392 460124 4396 460152
rect 4452 460124 4462 460180
rect 467954 459228 467964 459284
rect 468020 459228 469868 459284
rect 469924 459228 470120 459284
rect 12562 457772 12572 457828
rect 12628 457772 180684 457828
rect 180740 457772 180750 457828
rect 595560 456484 597000 456680
rect 590594 456428 590604 456484
rect 590660 456456 597000 456484
rect 590660 456428 595672 456456
rect 554428 455252 554484 455672
rect 554418 455196 554428 455252
rect 554484 455196 554494 455252
rect 467842 453180 467852 453236
rect 467908 453208 470680 453236
rect 467908 453180 470708 453208
rect 207554 452844 207564 452900
rect 207620 452844 246876 452900
rect 246932 452844 246942 452900
rect 4274 452732 4284 452788
rect 4340 452732 293132 452788
rect 293188 452732 293198 452788
rect 470652 452452 470708 453180
rect 470642 452396 470652 452452
rect 470708 452396 470718 452452
rect 470306 451500 470316 451556
rect 470372 451500 533036 451556
rect 533092 451500 533102 451556
rect 481618 451388 481628 451444
rect 481684 451388 558124 451444
rect 558180 451388 558190 451444
rect 481394 451276 481404 451332
rect 481460 451276 557788 451332
rect 557844 451276 557854 451332
rect 481506 451164 481516 451220
rect 481572 451164 557900 451220
rect 557956 451164 557966 451220
rect 187730 451052 187740 451108
rect 187796 451052 215740 451108
rect 215796 451052 215806 451108
rect 481282 451052 481292 451108
rect 481348 451052 558236 451108
rect 558292 451052 558302 451108
rect 478258 450604 478268 450660
rect 478324 450604 590828 450660
rect 590884 450604 590894 450660
rect 474870 450492 474908 450548
rect 474964 450492 474974 450548
rect 478482 450492 478492 450548
rect 478548 450492 590492 450548
rect 590548 450492 590558 450548
rect 467730 450380 467740 450436
rect 467796 450380 470876 450436
rect 470932 450380 470942 450436
rect 480498 450380 480508 450436
rect 480564 450380 554428 450436
rect 554484 450380 554494 450436
rect 468626 450268 468636 450324
rect 468692 450268 472892 450324
rect 472948 450268 472958 450324
rect 480610 450268 480620 450324
rect 480676 450268 558012 450324
rect 558068 450268 558078 450324
rect 532998 450156 533036 450212
rect 533092 450156 533102 450212
rect 459554 449596 459564 449652
rect 459620 449596 488124 449652
rect 488180 449596 488190 449652
rect 451266 449484 451276 449540
rect 451332 449484 504252 449540
rect 504308 449484 504318 449540
rect 7522 449372 7532 449428
rect 7588 449372 171724 449428
rect 171780 449372 171790 449428
rect 174290 449372 174300 449428
rect 174356 449372 218540 449428
rect 218596 449372 218606 449428
rect 449698 449372 449708 449428
rect 449764 449372 527436 449428
rect 527492 449372 527502 449428
rect 459442 448476 459452 448532
rect 459508 448476 521612 448532
rect 521668 448476 521678 448532
rect 526642 448476 526652 448532
rect 526708 448476 527436 448532
rect 527492 448476 531132 448532
rect 531188 448476 531198 448532
rect 474898 448364 474908 448420
rect 474964 448364 479612 448420
rect 479668 448364 479678 448420
rect 477922 447916 477932 447972
rect 477988 447916 493500 447972
rect 493556 447916 493566 447972
rect 478482 447804 478492 447860
rect 478548 447804 502908 447860
rect 502964 447804 502974 447860
rect 525746 447804 525756 447860
rect 525812 447804 540540 447860
rect 540596 447804 540606 447860
rect 475122 447692 475132 447748
rect 475188 447692 512316 447748
rect 512372 447692 512382 447748
rect 527090 447692 527100 447748
rect 527156 447692 549948 447748
rect 550004 447692 550014 447748
rect 521574 447356 521612 447412
rect 521668 447356 521678 447412
rect 480610 446908 480620 446964
rect 480676 446908 484092 446964
rect 484148 446908 484158 446964
rect 468626 446796 468636 446852
rect 468692 446796 474572 446852
rect 474628 446796 474638 446852
rect -960 446068 480 446264
rect 451042 446124 451052 446180
rect 451108 446124 509628 446180
rect 509684 446124 509694 446180
rect -960 446040 4956 446068
rect 392 446012 4956 446040
rect 5012 446012 5022 446068
rect 19282 446012 19292 446068
rect 19348 446012 167244 446068
rect 167300 446012 167310 446068
rect 452834 446012 452844 446068
rect 452900 446012 532700 446068
rect 532756 446012 532766 446068
rect 464482 444444 464492 444500
rect 464548 444444 482748 444500
rect 482804 444444 482814 444500
rect 152786 444332 152796 444388
rect 152852 444332 202412 444388
rect 202468 444332 202478 444388
rect 456194 444332 456204 444388
rect 456260 444332 506940 444388
rect 506996 444332 507006 444388
rect 595560 443268 597000 443464
rect 478034 443212 478044 443268
rect 478100 443240 597000 443268
rect 478100 443212 595672 443240
rect 190418 439292 190428 439348
rect 190484 439292 216748 439348
rect 216804 439292 216814 439348
rect 454514 439292 454524 439348
rect 454580 439292 532588 439348
rect 532644 439292 532654 439348
rect 185042 437948 185052 438004
rect 185108 437948 218428 438004
rect 218484 437948 218494 438004
rect 158162 437836 158172 437892
rect 158228 437836 214396 437892
rect 214452 437836 214462 437892
rect 456082 437836 456092 437892
rect 456148 437836 489468 437892
rect 489524 437836 489534 437892
rect 131282 437724 131292 437780
rect 131348 437724 214508 437780
rect 214564 437724 214574 437780
rect 457762 437724 457772 437780
rect 457828 437724 508284 437780
rect 508340 437724 508350 437780
rect 101714 437612 101724 437668
rect 101780 437612 288092 437668
rect 288148 437612 288158 437668
rect 451154 437612 451164 437668
rect 451220 437612 532812 437668
rect 532868 437612 532878 437668
rect 4386 436156 4396 436212
rect 4452 436156 298396 436212
rect 298452 436156 298462 436212
rect 4946 436044 4956 436100
rect 5012 436044 298844 436100
rect 298900 436044 298910 436100
rect 4162 435932 4172 435988
rect 4228 435932 298620 435988
rect 298676 435932 298686 435988
rect 142034 434476 142044 434532
rect 142100 434476 216860 434532
rect 216916 434476 216926 434532
rect 139346 434364 139356 434420
rect 139412 434364 216972 434420
rect 217028 434364 217038 434420
rect 449362 434364 449372 434420
rect 449428 434364 505596 434420
rect 505652 434364 505662 434420
rect 99026 434252 99036 434308
rect 99092 434252 279804 434308
rect 279860 434252 279870 434308
rect 452722 434252 452732 434308
rect 452788 434252 510972 434308
rect 511028 434252 511038 434308
rect 123218 433580 123228 433636
rect 123284 433580 295036 433636
rect 295092 433580 295102 433636
rect 117842 433468 117852 433524
rect 117908 433468 295260 433524
rect 295316 433468 295326 433524
rect 163538 433356 163548 433412
rect 163604 433356 164556 433412
rect 164612 433356 164622 433412
rect 166198 433356 166236 433412
rect 166292 433356 166302 433412
rect 169558 433356 169596 433412
rect 169652 433356 169662 433412
rect 265682 433356 265692 433412
rect 265748 433356 267036 433412
rect 267092 433356 267102 433412
rect 268678 433356 268716 433412
rect 268772 433356 268782 433412
rect 90962 432908 90972 432964
rect 91028 432908 300748 432964
rect 300804 432908 300814 432964
rect 464594 432908 464604 432964
rect 464660 432908 485436 432964
rect 485492 432908 485502 432964
rect 462802 432796 462812 432852
rect 462868 432796 484092 432852
rect 484148 432796 484158 432852
rect 107090 432684 107100 432740
rect 107156 432684 121772 432740
rect 121828 432684 121838 432740
rect 212482 432684 212492 432740
rect 212548 432684 272636 432740
rect 272692 432684 272702 432740
rect 461234 432684 461244 432740
rect 461300 432684 486780 432740
rect 486836 432684 486846 432740
rect 96338 432572 96348 432628
rect 96404 432572 121996 432628
rect 122052 432572 122062 432628
rect 209234 432572 209244 432628
rect 209300 432572 272972 432628
rect 273028 432572 273038 432628
rect 457762 432572 457772 432628
rect 457828 432572 490812 432628
rect 490868 432572 490878 432628
rect 512278 432572 512316 432628
rect 512372 432572 512382 432628
rect 206546 432460 206556 432516
rect 206612 432460 274764 432516
rect 274820 432460 274830 432516
rect 128594 432348 128604 432404
rect 128660 432348 298284 432404
rect 298340 432348 298350 432404
rect 112466 432236 112476 432292
rect 112532 432236 284844 432292
rect 284900 432236 284910 432292
rect 474562 432236 474572 432292
rect 474628 432236 497532 432292
rect 497588 432236 497598 432292
rect -960 431956 480 432152
rect 51986 432124 51996 432180
rect 52052 432124 66780 432180
rect 66836 432124 66846 432180
rect 115154 432124 115164 432180
rect 115220 432124 295148 432180
rect 295204 432124 295214 432180
rect 482962 432124 482972 432180
rect 483028 432124 496188 432180
rect 496244 432124 496254 432180
rect 498838 432124 498876 432180
rect 498932 432124 498942 432180
rect 64082 432012 64092 432068
rect 64148 432012 76412 432068
rect 76468 432012 76478 432068
rect 88274 432012 88284 432068
rect 88340 432012 276444 432068
rect 276500 432012 276510 432068
rect 478370 432012 478380 432068
rect 478436 432012 492156 432068
rect 492212 432012 492222 432068
rect 502870 432012 502908 432068
rect 502964 432012 502974 432068
rect -960 431928 4956 431956
rect 392 431900 4956 431928
rect 5012 431900 5022 431956
rect 60386 431900 60396 431956
rect 60452 431900 72156 431956
rect 72212 431900 72222 431956
rect 82870 431900 82908 431956
rect 82964 431900 82974 431956
rect 85586 431900 85596 431956
rect 85652 431900 279804 431956
rect 279860 431900 279870 431956
rect 478146 431900 478156 431956
rect 478212 431900 494844 431956
rect 494900 431900 494910 431956
rect 518998 431900 519036 431956
rect 519092 431900 519102 431956
rect 77494 431788 77532 431844
rect 77588 431788 77598 431844
rect 483074 431788 483084 431844
rect 483140 431788 493500 431844
rect 493556 431788 493566 431844
rect 523030 431788 523068 431844
rect 523124 431788 523134 431844
rect 257618 431004 257628 431060
rect 257684 431004 300860 431060
rect 300916 431004 300926 431060
rect 254930 430892 254940 430948
rect 254996 430892 301084 430948
rect 301140 430892 301150 430948
rect 244178 430780 244188 430836
rect 244244 430780 301084 430836
rect 301140 430780 301150 430836
rect 219986 430668 219996 430724
rect 220052 430668 288092 430724
rect 288148 430668 288158 430724
rect 203858 430556 203868 430612
rect 203924 430556 278012 430612
rect 278068 430556 278078 430612
rect 214610 430444 214620 430500
rect 214676 430444 298284 430500
rect 298340 430444 298350 430500
rect 55234 430332 55244 430388
rect 55300 430332 193116 430388
rect 193172 430332 193182 430388
rect 201170 430332 201180 430388
rect 201236 430332 293244 430388
rect 293300 430332 293310 430388
rect 69430 430220 69468 430276
rect 69524 430220 69534 430276
rect 93650 430220 93660 430276
rect 93716 430220 298620 430276
rect 298676 430220 298686 430276
rect 464594 430220 464604 430276
rect 464660 430220 521724 430276
rect 521780 430220 521790 430276
rect 595560 430164 597000 430248
rect 56914 430108 56924 430164
rect 56980 430108 294924 430164
rect 294980 430108 294990 430164
rect 462802 430108 462812 430164
rect 462868 430108 524412 430164
rect 524468 430108 524478 430164
rect 590818 430108 590828 430164
rect 590884 430108 597000 430164
rect 66658 429996 66668 430052
rect 66724 429996 212492 430052
rect 212548 429996 212558 430052
rect 212818 429996 212828 430052
rect 212884 429996 278124 430052
rect 278180 429996 278190 430052
rect 456082 429996 456092 430052
rect 456148 429996 519596 430052
rect 519652 429996 519662 430052
rect 595560 430024 597000 430108
rect 56466 429884 56476 429940
rect 56532 429884 300972 429940
rect 301028 429884 301038 429940
rect 478370 429884 478380 429940
rect 478436 429884 513660 429940
rect 513716 429884 513726 429940
rect 4610 429772 4620 429828
rect 4676 429772 298060 429828
rect 298116 429772 298126 429828
rect 477586 429772 477596 429828
rect 477652 429772 515004 429828
rect 515060 429772 515070 429828
rect 4386 429660 4396 429716
rect 4452 429660 298508 429716
rect 298564 429660 298574 429716
rect 477810 429660 477820 429716
rect 477876 429660 516348 429716
rect 516404 429660 516414 429716
rect 4162 429548 4172 429604
rect 4228 429548 298732 429604
rect 298788 429548 298798 429604
rect 449474 429548 449484 429604
rect 449540 429548 532924 429604
rect 532980 429548 532990 429604
rect 80210 429436 80220 429492
rect 80276 429436 291564 429492
rect 291620 429436 291630 429492
rect 478146 429436 478156 429492
rect 478212 429436 517692 429492
rect 517748 429436 517758 429492
rect 74806 429324 74844 429380
rect 74900 429324 74910 429380
rect 196532 429324 231868 429380
rect 196532 429268 196588 429324
rect 231812 429268 231868 429324
rect 243572 429324 267148 429380
rect 461122 429324 461132 429380
rect 461188 429324 500220 429380
rect 500276 429324 500286 429380
rect 243572 429268 243628 429324
rect 267092 429268 267148 429324
rect 125906 429212 125916 429268
rect 125972 429212 196588 429268
rect 217298 429212 217308 429268
rect 217364 429212 220108 429268
rect 231812 429212 243628 429268
rect 249526 429212 249564 429268
rect 249620 429212 249630 429268
rect 252214 429212 252252 429268
rect 252308 429212 252318 429268
rect 260278 429212 260316 429268
rect 260372 429212 260382 429268
rect 262994 429212 263004 429268
rect 263060 429212 263676 429268
rect 263732 429212 263742 429268
rect 267092 429212 289884 429268
rect 289940 429212 289950 429268
rect 464482 429212 464492 429268
rect 464548 429212 501564 429268
rect 501620 429212 501630 429268
rect 220052 429156 220108 429212
rect 220052 429100 279692 429156
rect 279748 429100 279758 429156
rect 60582 428540 60620 428596
rect 60676 428540 60686 428596
rect 83234 428428 83244 428484
rect 83300 428428 298956 428484
rect 299012 428428 299022 428484
rect 252242 427756 252252 427812
rect 252308 427756 301084 427812
rect 301140 427756 301150 427812
rect 249554 427644 249564 427700
rect 249620 427644 300860 427700
rect 300916 427644 300926 427700
rect 83570 427532 83580 427588
rect 83636 427532 295260 427588
rect 295316 427532 295326 427588
rect 83346 427420 83356 427476
rect 83412 427420 295036 427476
rect 295092 427420 295102 427476
rect 56802 427308 56812 427364
rect 56868 427308 284956 427364
rect 285012 427308 285022 427364
rect 56690 427196 56700 427252
rect 56756 427196 296492 427252
rect 296548 427196 296558 427252
rect 56354 427084 56364 427140
rect 56420 427084 300860 427140
rect 300916 427084 300926 427140
rect 480060 426916 480116 427560
rect 480050 426860 480060 426916
rect 480116 426860 480126 426916
rect 529928 426412 532588 426468
rect 532644 426412 532654 426468
rect 478706 425964 478716 426020
rect 478772 425964 480088 426020
rect 60060 425124 60116 425768
rect 60050 425068 60060 425124
rect 60116 425068 60126 425124
rect 60172 423892 60228 424424
rect 478594 424396 478604 424452
rect 478660 424396 480088 424452
rect 60162 423836 60172 423892
rect 60228 423836 60238 423892
rect 58370 423052 58380 423108
rect 58436 423052 60088 423108
rect 477026 422828 477036 422884
rect 477092 422828 480088 422884
rect 269864 422380 270620 422436
rect 270676 422380 270686 422436
rect 60284 421652 60340 421736
rect 60274 421596 60284 421652
rect 60340 421596 60350 421652
rect 468626 421260 468636 421316
rect 468692 421260 480088 421316
rect 269864 421036 270732 421092
rect 270788 421036 270798 421092
rect 529928 421036 532700 421092
rect 532756 421036 532766 421092
rect 50194 420364 50204 420420
rect 50260 420364 60088 420420
rect 269864 419692 270844 419748
rect 270900 419692 270910 419748
rect 476914 419692 476924 419748
rect 476980 419692 480088 419748
rect 58258 419020 58268 419076
rect 58324 419020 60088 419076
rect 269864 418348 273980 418404
rect 274036 418348 274046 418404
rect 460226 418124 460236 418180
rect 460292 418124 480088 418180
rect 392 418040 4620 418068
rect -960 418012 4620 418040
rect 4676 418012 4686 418068
rect -960 417816 480 418012
rect 58146 417676 58156 417732
rect 58212 417676 60088 417732
rect 269864 417004 275548 417060
rect 275604 417004 275614 417060
rect 595560 416836 597000 417032
rect 590706 416780 590716 416836
rect 590772 416808 597000 416836
rect 590772 416780 595672 416808
rect 460114 416556 460124 416612
rect 460180 416556 480088 416612
rect 48626 416332 48636 416388
rect 48692 416332 60088 416388
rect 269864 415660 273868 415716
rect 273924 415660 273934 415716
rect 529928 415660 532812 415716
rect 532868 415660 532878 415716
rect 49970 414988 49980 415044
rect 50036 414988 60088 415044
rect 476242 414988 476252 415044
rect 476308 414988 480088 415044
rect 269864 414316 272188 414372
rect 272244 414316 272254 414372
rect 56578 413644 56588 413700
rect 56644 413644 60088 413700
rect 476466 413420 476476 413476
rect 476532 413420 480088 413476
rect 269864 412972 272300 413028
rect 272356 412972 272366 413028
rect 57026 412300 57036 412356
rect 57092 412300 60088 412356
rect 451042 411852 451052 411908
rect 451108 411852 480088 411908
rect 269864 411628 272412 411684
rect 272468 411628 272478 411684
rect 56690 410956 56700 411012
rect 56756 410956 60088 411012
rect 269500 410004 269556 410312
rect 449362 410284 449372 410340
rect 449428 410284 480088 410340
rect 529928 410284 532924 410340
rect 532980 410284 532990 410340
rect 269490 409948 269500 410004
rect 269556 409948 269566 410004
rect 56802 409612 56812 409668
rect 56868 409612 60088 409668
rect 60162 409164 60172 409220
rect 60228 409164 60238 409220
rect 60172 408296 60228 409164
rect 269864 408940 270508 408996
rect 270564 408940 270574 408996
rect 456082 408716 456092 408772
rect 456148 408716 480088 408772
rect 60274 407708 60284 407764
rect 60340 407708 60350 407764
rect 60284 406952 60340 407708
rect 269864 407596 272524 407652
rect 272580 407596 272590 407652
rect 533362 407372 533372 407428
rect 533428 407372 554428 407428
rect 554484 407372 554494 407428
rect 452722 407148 452732 407204
rect 452788 407148 480088 407204
rect 269388 405748 269444 406280
rect 269378 405692 269388 405748
rect 269444 405692 269454 405748
rect 56914 405580 56924 405636
rect 56980 405580 60088 405636
rect 474786 405580 474796 405636
rect 474852 405580 480088 405636
rect 269864 404908 270956 404964
rect 271012 404908 271022 404964
rect 529928 404908 533372 404964
rect 533428 404908 533438 404964
rect 60396 404684 60508 404740
rect 60564 404684 60574 404740
rect 60396 404264 60452 404684
rect 454402 404012 454412 404068
rect 454468 404012 480088 404068
rect 392 403928 4284 403956
rect -960 403900 4284 403928
rect 4340 403900 4350 403956
rect -960 403704 480 403900
rect 595560 403620 597000 403816
rect 269864 403564 275660 403620
rect 275716 403564 275726 403620
rect 591042 403564 591052 403620
rect 591108 403592 597000 403620
rect 591108 403564 595672 403592
rect 468626 403340 468636 403396
rect 468692 403340 469980 403396
rect 470036 403340 470046 403396
rect 478772 403116 480620 403172
rect 480676 403116 480686 403172
rect 50082 402892 50092 402948
rect 50148 402892 60088 402948
rect 284722 402892 284732 402948
rect 284788 402892 476252 402948
rect 476308 402892 476318 402948
rect 288082 402780 288092 402836
rect 288148 402780 476476 402836
rect 476532 402780 476542 402836
rect 478772 402724 478828 403116
rect 301746 402668 301756 402724
rect 301812 402668 478828 402724
rect 298610 402556 298620 402612
rect 298676 402556 478380 402612
rect 478436 402556 478446 402612
rect 472882 402444 472892 402500
rect 472948 402444 480088 402500
rect 300738 402332 300748 402388
rect 300804 402332 478044 402388
rect 478100 402332 478110 402388
rect 269864 402220 274092 402276
rect 274148 402220 274158 402276
rect 298834 402220 298844 402276
rect 298900 402220 477596 402276
rect 477652 402220 477662 402276
rect 48402 401548 48412 401604
rect 48468 401548 60088 401604
rect 295138 401436 295148 401492
rect 295204 401436 477932 401492
rect 477988 401436 477998 401492
rect 298050 401324 298060 401380
rect 298116 401324 478156 401380
rect 478212 401324 478222 401380
rect 298386 401212 298396 401268
rect 298452 401212 478380 401268
rect 478436 401212 478446 401268
rect 300850 401100 300860 401156
rect 300916 401100 480508 401156
rect 480564 401100 480574 401156
rect 269864 400876 278124 400932
rect 278180 400876 278190 400932
rect 474674 400876 474684 400932
rect 474740 400876 480088 400932
rect 301634 400652 301644 400708
rect 301700 400652 480508 400708
rect 480564 400652 480574 400708
rect 301522 400540 301532 400596
rect 301588 400540 480620 400596
rect 480676 400540 480686 400596
rect 301074 400428 301084 400484
rect 301140 400428 455308 400484
rect 455252 400260 455308 400428
rect 56914 400204 56924 400260
rect 56980 400204 60088 400260
rect 455252 400204 480620 400260
rect 480676 400204 480686 400260
rect 295250 399756 295260 399812
rect 295316 399756 478492 399812
rect 478548 399756 478558 399812
rect 298050 399644 298060 399700
rect 298116 399644 477820 399700
rect 477876 399644 477886 399700
rect 269864 399532 291452 399588
rect 291508 399532 291518 399588
rect 298498 399532 298508 399588
rect 298564 399532 478044 399588
rect 478100 399532 478110 399588
rect 529928 399532 549500 399588
rect 549556 399532 549566 399588
rect 298946 399420 298956 399476
rect 299012 399420 478268 399476
rect 478324 399420 478334 399476
rect 474562 399308 474572 399364
rect 474628 399308 480088 399364
rect 51762 398860 51772 398916
rect 51828 398860 60088 398916
rect 269864 398188 274652 398244
rect 274708 398188 274718 398244
rect 295026 398076 295036 398132
rect 295092 398076 475132 398132
rect 475188 398076 475198 398132
rect 298162 397964 298172 398020
rect 298228 397964 478156 398020
rect 478212 397964 478222 398020
rect 468514 397740 468524 397796
rect 468580 397740 480088 397796
rect 48514 397516 48524 397572
rect 48580 397516 60088 397572
rect 272962 397292 272972 397348
rect 273028 397292 476252 397348
rect 476308 397292 476318 397348
rect 269864 396844 293132 396900
rect 293188 396844 293198 396900
rect 56690 396172 56700 396228
rect 56756 396172 60088 396228
rect 468402 396172 468412 396228
rect 468468 396172 480088 396228
rect 269864 395500 299852 395556
rect 299908 395500 299918 395556
rect 56242 394828 56252 394884
rect 56308 394828 60088 394884
rect 468290 394604 468300 394660
rect 468356 394604 480088 394660
rect 269864 394156 294812 394212
rect 294868 394156 294878 394212
rect 529928 394156 549388 394212
rect 549444 394156 549454 394212
rect 56802 393484 56812 393540
rect 56868 393484 60088 393540
rect 468178 393036 468188 393092
rect 468244 393036 480088 393092
rect 269864 392812 296492 392868
rect 296548 392812 296558 392868
rect 56690 392140 56700 392196
rect 56756 392140 60088 392196
rect 269864 391468 298172 391524
rect 298228 391468 298238 391524
rect 470082 391468 470092 391524
rect 470148 391468 480088 391524
rect 56802 390796 56812 390852
rect 56868 390796 60088 390852
rect 273186 390572 273196 390628
rect 273252 390572 474796 390628
rect 474852 390572 474862 390628
rect 533362 390572 533372 390628
rect 533428 390572 548156 390628
rect 548212 390572 548222 390628
rect 595560 390404 597000 390600
rect 590930 390348 590940 390404
rect 590996 390376 597000 390404
rect 590996 390348 595672 390376
rect 269864 390124 289772 390180
rect 289828 390124 289838 390180
rect 470866 389900 470876 389956
rect 470932 389900 480088 389956
rect -960 389732 480 389816
rect -960 389676 4396 389732
rect 4452 389676 4462 389732
rect -960 389592 480 389676
rect 56466 389452 56476 389508
rect 56532 389452 60088 389508
rect 269864 388780 272636 388836
rect 272692 388780 273532 388836
rect 273588 388780 273598 388836
rect 529928 388780 533372 388836
rect 533428 388780 533438 388836
rect 472882 388332 472892 388388
rect 472948 388332 480088 388388
rect 56914 388108 56924 388164
rect 56980 388108 60088 388164
rect 269864 387436 451052 387492
rect 451108 387436 451118 387492
rect 56354 386764 56364 386820
rect 56420 386764 60088 386820
rect 469970 386764 469980 386820
rect 470036 386764 480088 386820
rect 269864 386092 449372 386148
rect 449428 386092 449438 386148
rect 56130 385420 56140 385476
rect 56196 385420 60088 385476
rect 470194 385196 470204 385252
rect 470260 385196 480088 385252
rect 269864 384748 456092 384804
rect 456148 384748 456158 384804
rect 60284 383348 60340 384104
rect 273634 383964 273644 384020
rect 273700 383964 472892 384020
rect 472948 383964 472958 384020
rect 274754 383852 274764 383908
rect 274820 383852 476364 383908
rect 476420 383852 476430 383908
rect 469858 383628 469868 383684
rect 469924 383628 480088 383684
rect 269864 383404 452732 383460
rect 452788 383404 452798 383460
rect 529928 383404 533036 383460
rect 533092 383404 533102 383460
rect 60274 383292 60284 383348
rect 60340 383292 60350 383348
rect 53666 382732 53676 382788
rect 53732 382732 60088 382788
rect 269864 382060 273196 382116
rect 273252 382060 273262 382116
rect 470642 382060 470652 382116
rect 470708 382060 480088 382116
rect 279682 381836 279692 381892
rect 279748 381836 484764 381892
rect 484820 381836 484830 381892
rect 54338 381388 54348 381444
rect 54404 381388 60088 381444
rect 272962 381388 272972 381444
rect 273028 381388 459452 381444
rect 459508 381388 459518 381444
rect 269864 380716 454412 380772
rect 454468 380716 454478 380772
rect 484726 380716 484764 380772
rect 484820 380716 484830 380772
rect 273746 380604 273756 380660
rect 273812 380604 474684 380660
rect 474740 380604 474750 380660
rect 502292 380604 525868 380660
rect 502292 380548 502348 380604
rect 279794 380492 279804 380548
rect 279860 380492 502348 380548
rect 525812 380548 525868 380604
rect 525812 380492 590604 380548
rect 590660 380492 590670 380548
rect 300962 380380 300972 380436
rect 301028 380380 502908 380436
rect 502964 380380 502974 380436
rect 525858 380380 525868 380436
rect 525924 380380 526316 380436
rect 526372 380380 526382 380436
rect 298498 380268 298508 380324
rect 298564 380268 500892 380324
rect 500948 380268 500958 380324
rect 278002 380156 278012 380212
rect 278068 380156 482748 380212
rect 482804 380156 482814 380212
rect 490532 380156 502348 380212
rect 490532 380100 490588 380156
rect 502292 380100 502348 380156
rect 57922 380044 57932 380100
rect 57988 380044 60088 380100
rect 298274 380044 298284 380100
rect 298340 380044 490588 380100
rect 492818 380044 492828 380100
rect 492884 380044 492894 380100
rect 502292 380044 523068 380100
rect 523124 380044 523134 380100
rect 492828 379988 492884 380044
rect 459442 379932 459452 379988
rect 459508 379932 492884 379988
rect 284834 379596 284844 379652
rect 284900 379596 519036 379652
rect 519092 379596 519102 379652
rect 294914 379484 294924 379540
rect 294980 379484 496860 379540
rect 496916 379484 496926 379540
rect 269864 379372 273644 379428
rect 273700 379372 273710 379428
rect 479602 379372 479612 379428
rect 479668 379372 515004 379428
rect 515060 379372 515070 379428
rect 476914 379036 476924 379092
rect 476980 379036 559468 379092
rect 559524 379036 559534 379092
rect 299058 378924 299068 378980
rect 299124 378924 517020 378980
rect 517076 378924 517086 378980
rect 276322 378812 276332 378868
rect 276388 378812 590492 378868
rect 590548 378812 590558 378868
rect 53554 378700 53564 378756
rect 53620 378700 60088 378756
rect 269864 378028 273756 378084
rect 273812 378028 273822 378084
rect 494806 377916 494844 377972
rect 494900 377916 494910 377972
rect 498838 377916 498876 377972
rect 498932 377916 498942 377972
rect 521014 377916 521052 377972
rect 521108 377916 521118 377972
rect 521602 377916 521612 377972
rect 521668 377916 525084 377972
rect 525140 377916 525150 377972
rect 461122 377804 461132 377860
rect 461188 377804 488796 377860
rect 488852 377804 488862 377860
rect 462914 377692 462924 377748
rect 462980 377692 486780 377748
rect 486836 377692 486846 377748
rect 454402 377580 454412 377636
rect 454468 377580 490812 377636
rect 490868 377580 490878 377636
rect 478146 377468 478156 377524
rect 478212 377468 504924 377524
rect 504980 377468 504990 377524
rect 56802 377356 56812 377412
rect 56868 377356 60088 377412
rect 477922 377356 477932 377412
rect 477988 377356 508956 377412
rect 509012 377356 509022 377412
rect 479602 377244 479612 377300
rect 479668 377244 510972 377300
rect 511028 377244 511038 377300
rect 595560 377188 597000 377384
rect 467842 377132 467852 377188
rect 467908 377132 512988 377188
rect 513044 377132 513054 377188
rect 590146 377132 590156 377188
rect 590212 377160 597000 377188
rect 590212 377132 595672 377160
rect 269864 376684 299068 376740
rect 299124 376684 299134 376740
rect 392 375704 4172 375732
rect -960 375676 4172 375704
rect 4228 375676 4238 375732
rect -960 375480 480 375676
rect 60172 375396 60228 376040
rect 477026 375452 477036 375508
rect 477092 375452 559580 375508
rect 559636 375452 559646 375508
rect 60162 375340 60172 375396
rect 60228 375340 60238 375396
rect 269864 375340 294924 375396
rect 294980 375340 294990 375396
rect 60722 374668 60732 374724
rect 60788 374668 60798 374724
rect 269864 373996 289772 374052
rect 289828 373996 289838 374052
rect 478594 373772 478604 373828
rect 478660 373772 563500 373828
rect 563556 373772 563566 373828
rect 56690 373324 56700 373380
rect 56756 373324 60088 373380
rect 269864 372652 296492 372708
rect 296548 372652 296558 372708
rect 478706 372092 478716 372148
rect 478772 372092 569212 372148
rect 569268 372092 569278 372148
rect 56578 371980 56588 372036
rect 56644 371980 60088 372036
rect 269864 371308 273756 371364
rect 273812 371308 273822 371364
rect 269864 369964 272972 370020
rect 273028 369964 273038 370020
rect 60172 368676 60228 369320
rect 480050 368844 480060 368900
rect 480116 368844 574924 368900
rect 574980 368844 574990 368900
rect 388882 368732 388892 368788
rect 388948 368732 506940 368788
rect 506996 368732 507006 368788
rect 60162 368620 60172 368676
rect 60228 368620 60238 368676
rect 269864 368620 273756 368676
rect 273812 368620 273822 368676
rect 60722 367948 60732 368004
rect 60788 367948 60798 368004
rect 269864 367276 273756 367332
rect 273812 367276 273822 367332
rect 60722 366604 60732 366660
rect 60788 366604 60798 366660
rect 269864 365932 273756 365988
rect 273812 365932 273822 365988
rect 58482 365260 58492 365316
rect 58548 365260 60088 365316
rect 269864 364588 273756 364644
rect 273812 364588 273822 364644
rect 590594 364140 590604 364196
rect 590660 364168 595672 364196
rect 590660 364140 597000 364168
rect 60050 363916 60060 363972
rect 60116 363916 60126 363972
rect 595560 363944 597000 364140
rect 269864 363244 273084 363300
rect 273140 363244 273150 363300
rect 56466 362572 56476 362628
rect 56532 362572 60088 362628
rect 269864 361900 273756 361956
rect 273812 361900 273822 361956
rect 392 361592 4172 361620
rect -960 361564 4172 361592
rect 4228 361564 4238 361620
rect -960 361368 480 361564
rect 55010 361228 55020 361284
rect 55076 361228 60088 361284
rect 269864 360556 273756 360612
rect 273812 360556 273822 360612
rect 56354 359884 56364 359940
rect 56420 359884 60088 359940
rect 269864 359212 273308 359268
rect 273364 359212 273374 359268
rect 54786 358540 54796 358596
rect 54852 358540 60088 358596
rect 269864 357868 273644 357924
rect 273700 357868 273710 357924
rect 53442 357196 53452 357252
rect 53508 357196 60088 357252
rect 269864 356524 273756 356580
rect 273812 356524 273822 356580
rect 53218 355852 53228 355908
rect 53284 355852 60088 355908
rect 269864 355180 273756 355236
rect 273812 355180 273822 355236
rect 53330 354508 53340 354564
rect 53396 354508 60088 354564
rect 56690 354396 56700 354452
rect 56756 354396 59612 354452
rect 59668 354396 59678 354452
rect 269864 353836 299852 353892
rect 299908 353836 299918 353892
rect 56242 353164 56252 353220
rect 56308 353164 60088 353220
rect 269864 352492 294812 352548
rect 294868 352492 294878 352548
rect 54898 351820 54908 351876
rect 54964 351820 60088 351876
rect 269864 351148 273644 351204
rect 273700 351148 273710 351204
rect 595560 350756 597000 350952
rect 591042 350700 591052 350756
rect 591108 350728 597000 350756
rect 591108 350700 595672 350728
rect 60396 350084 60452 350504
rect 60396 350028 60508 350084
rect 60564 350028 60574 350084
rect 269864 349804 273756 349860
rect 273812 349804 273822 349860
rect 54674 349132 54684 349188
rect 54740 349132 60088 349188
rect 482514 348572 482524 348628
rect 482580 348572 521612 348628
rect 521668 348572 521678 348628
rect 269864 348460 273756 348516
rect 273812 348460 273822 348516
rect 54562 347788 54572 347844
rect 54628 347788 60088 347844
rect 269602 347788 269612 347844
rect 269668 347788 272524 347844
rect 272580 347788 272590 347844
rect 392 347480 4172 347508
rect -960 347452 4172 347480
rect 4228 347452 4238 347508
rect -960 347256 480 347452
rect 269864 347116 284732 347172
rect 284788 347116 284798 347172
rect 60274 346444 60284 346500
rect 60340 346444 60350 346500
rect 269864 345772 291452 345828
rect 291508 345772 291518 345828
rect 498950 345324 498988 345380
rect 499044 345324 499054 345380
rect 502338 345324 502348 345380
rect 502404 345324 502442 345380
rect 505670 345324 505708 345380
rect 505764 345324 505774 345380
rect 60396 344484 60452 345128
rect 495926 344876 495964 344932
rect 496020 344876 496030 344932
rect 479938 344652 479948 344708
rect 480004 344652 492604 344708
rect 492660 344652 492670 344708
rect 479714 344540 479724 344596
rect 479780 344540 485884 344596
rect 485940 344540 485950 344596
rect 60396 344428 60508 344484
rect 60564 344428 60574 344484
rect 269864 344428 272972 344484
rect 273028 344428 273038 344484
rect 480162 344428 480172 344484
rect 480228 344428 489244 344484
rect 489300 344428 489310 344484
rect 509366 344428 509404 344484
rect 509460 344428 509470 344484
rect 512726 344428 512764 344484
rect 512820 344428 512830 344484
rect 516086 344428 516124 344484
rect 516180 344428 516190 344484
rect 519446 344428 519484 344484
rect 519540 344428 519550 344484
rect 58482 343756 58492 343812
rect 58548 343756 60088 343812
rect 269864 343084 293132 343140
rect 293188 343084 293198 343140
rect 419122 342748 419132 342804
rect 419188 342748 482524 342804
rect 482580 342748 482590 342804
rect 50306 342412 50316 342468
rect 50372 342412 60088 342468
rect 269864 341740 273196 341796
rect 273252 341740 273262 341796
rect 55346 341068 55356 341124
rect 55412 341068 60088 341124
rect 269864 340396 273756 340452
rect 273812 340396 273822 340452
rect 53666 339724 53676 339780
rect 53732 339724 60088 339780
rect 269864 339052 298172 339108
rect 298228 339052 298238 339108
rect 51986 338380 51996 338436
rect 52052 338380 60088 338436
rect 475458 338380 475468 338436
rect 475524 338380 480088 338436
rect 269864 337708 273308 337764
rect 273364 337708 273374 337764
rect 595560 337540 597000 337736
rect 475458 337484 475468 337540
rect 475524 337484 480088 337540
rect 591154 337484 591164 337540
rect 591220 337512 597000 337540
rect 591220 337484 595672 337512
rect 58706 337036 58716 337092
rect 58772 337036 60088 337092
rect 475570 336588 475580 336644
rect 475636 336588 480088 336644
rect 269864 336364 273084 336420
rect 273140 336364 273150 336420
rect 60722 335692 60732 335748
rect 60788 335692 60798 335748
rect 475458 335692 475468 335748
rect 475524 335692 480088 335748
rect 60162 335020 60172 335076
rect 60228 335020 60238 335076
rect 269864 335020 273084 335076
rect 273140 335020 273150 335076
rect 60172 334376 60228 335020
rect 476242 334796 476252 334852
rect 476308 334796 480088 334852
rect 271282 334348 271292 334404
rect 271348 334348 272412 334404
rect 272468 334348 272478 334404
rect 476354 333900 476364 333956
rect 476420 333900 480088 333956
rect 269864 333676 272972 333732
rect 273028 333676 273038 333732
rect -960 333172 480 333368
rect -960 333144 4172 333172
rect 392 333116 4172 333144
rect 4228 333116 4238 333172
rect 60498 333004 60508 333060
rect 60564 333004 60574 333060
rect 475458 333004 475468 333060
rect 475524 333004 480088 333060
rect 269864 332332 273196 332388
rect 273252 332332 273262 332388
rect 475458 332108 475468 332164
rect 475524 332108 480088 332164
rect 53106 331660 53116 331716
rect 53172 331660 60088 331716
rect 475570 331212 475580 331268
rect 475636 331212 480088 331268
rect 269864 330988 284732 331044
rect 284788 330988 284798 331044
rect 60172 329476 60228 330344
rect 475458 330316 475468 330372
rect 475524 330316 480088 330372
rect 269864 329644 298172 329700
rect 298228 329644 298238 329700
rect 60162 329420 60172 329476
rect 60228 329420 60238 329476
rect 475682 329420 475692 329476
rect 475748 329420 480088 329476
rect 58146 328972 58156 329028
rect 58212 328972 60088 329028
rect 390562 328524 390572 328580
rect 390628 328524 480088 328580
rect 269864 328300 273308 328356
rect 273364 328300 273374 328356
rect 60722 327628 60732 327684
rect 60788 327628 60798 327684
rect 476242 327628 476252 327684
rect 476308 327628 480088 327684
rect 269864 326956 273532 327012
rect 273588 326956 273598 327012
rect 475458 326732 475468 326788
rect 475524 326732 480088 326788
rect 58258 326284 58268 326340
rect 58324 326284 60088 326340
rect 476466 325836 476476 325892
rect 476532 325836 480088 325892
rect 269864 325612 273420 325668
rect 273476 325612 273486 325668
rect 60396 324324 60452 324968
rect 476242 324940 476252 324996
rect 476308 324940 480088 324996
rect 590482 324492 590492 324548
rect 590548 324520 595672 324548
rect 590548 324492 597000 324520
rect 53666 324268 53676 324324
rect 53732 324268 56252 324324
rect 56308 324268 56318 324324
rect 60386 324268 60396 324324
rect 60452 324268 60462 324324
rect 269864 324268 293132 324324
rect 293188 324268 293198 324324
rect 595560 324296 597000 324492
rect 476690 324044 476700 324100
rect 476756 324044 480088 324100
rect 58034 323596 58044 323652
rect 58100 323596 60088 323652
rect 476914 323148 476924 323204
rect 476980 323148 480088 323204
rect 269864 322924 291452 322980
rect 291508 322924 291518 322980
rect 55234 322252 55244 322308
rect 55300 322252 60088 322308
rect 476354 322252 476364 322308
rect 476420 322252 480088 322308
rect 269864 321580 296492 321636
rect 296548 321580 296558 321636
rect 475458 321356 475468 321412
rect 475524 321356 480088 321412
rect 58370 320908 58380 320964
rect 58436 320908 60088 320964
rect 472882 320460 472892 320516
rect 472948 320460 480088 320516
rect 269864 320236 299852 320292
rect 299908 320236 299918 320292
rect 54450 319564 54460 319620
rect 54516 319564 60088 319620
rect 473106 319564 473116 319620
rect 473172 319564 480088 319620
rect -960 319060 480 319256
rect -960 319032 4284 319060
rect 392 319004 4284 319032
rect 4340 319004 4350 319060
rect 269864 318892 273756 318948
rect 273812 318892 273822 318948
rect 475570 318668 475580 318724
rect 475636 318668 480088 318724
rect 57026 318220 57036 318276
rect 57092 318220 60088 318276
rect 475458 317772 475468 317828
rect 475524 317772 480088 317828
rect 269864 317548 294812 317604
rect 294868 317548 294878 317604
rect 58594 316876 58604 316932
rect 58660 316876 60088 316932
rect 476802 316876 476812 316932
rect 476868 316876 480088 316932
rect 269864 316204 289772 316260
rect 289828 316204 289838 316260
rect 477026 315980 477036 316036
rect 477092 315980 480088 316036
rect 58706 315532 58716 315588
rect 58772 315532 60088 315588
rect 475458 315084 475468 315140
rect 475524 315084 480088 315140
rect 269864 314860 288092 314916
rect 288148 314860 288158 314916
rect 51874 314188 51884 314244
rect 51940 314188 60088 314244
rect 476578 314188 476588 314244
rect 476644 314188 480088 314244
rect 269864 313516 279692 313572
rect 279748 313516 279758 313572
rect 475458 313292 475468 313348
rect 475524 313292 480088 313348
rect 50306 312844 50316 312900
rect 50372 312844 60088 312900
rect 476130 312396 476140 312452
rect 476196 312396 480088 312452
rect 269864 312172 277676 312228
rect 277732 312172 277742 312228
rect 55346 311500 55356 311556
rect 55412 311500 60088 311556
rect 476578 311500 476588 311556
rect 476644 311500 480088 311556
rect 595560 311108 597000 311304
rect 591266 311052 591276 311108
rect 591332 311080 597000 311108
rect 591332 311052 595672 311080
rect 269864 310828 272188 310884
rect 272244 310828 272254 310884
rect 476914 310604 476924 310660
rect 476980 310604 480088 310660
rect 58706 310156 58716 310212
rect 58772 310156 60088 310212
rect 476354 309708 476364 309764
rect 476420 309708 480088 309764
rect 269864 309484 279020 309540
rect 279076 309484 279086 309540
rect 58594 308812 58604 308868
rect 58660 308812 60088 308868
rect 475458 308812 475468 308868
rect 475524 308812 480088 308868
rect 269864 308140 273868 308196
rect 273924 308140 273934 308196
rect 476242 307916 476252 307972
rect 476308 307916 480088 307972
rect 60722 307468 60732 307524
rect 60788 307468 60798 307524
rect 56802 307356 56812 307412
rect 56868 307356 59836 307412
rect 59892 307356 59902 307412
rect 476690 307020 476700 307076
rect 476756 307020 480088 307076
rect 269864 306796 278908 306852
rect 278964 306796 278974 306852
rect 269826 306236 269836 306292
rect 269892 306236 272300 306292
rect 272356 306236 272366 306292
rect 57026 306124 57036 306180
rect 57092 306124 60088 306180
rect 476466 306124 476476 306180
rect 476532 306124 480088 306180
rect 269864 305452 278796 305508
rect 278852 305452 278862 305508
rect 476130 305228 476140 305284
rect 476196 305228 480088 305284
rect -960 304948 480 305144
rect -960 304920 4396 304948
rect 392 304892 4396 304920
rect 4452 304892 4462 304948
rect 60274 304780 60284 304836
rect 60340 304780 60350 304836
rect 476802 304332 476812 304388
rect 476868 304332 480088 304388
rect 269724 304052 269780 304136
rect 269714 303996 269724 304052
rect 269780 303996 269790 304052
rect 55122 303436 55132 303492
rect 55188 303436 60088 303492
rect 477026 303436 477036 303492
rect 477092 303436 480088 303492
rect 269864 302764 272300 302820
rect 272356 302764 272366 302820
rect 388098 302316 388108 302372
rect 388164 302316 476924 302372
rect 476980 302316 476990 302372
rect 56018 302092 56028 302148
rect 56084 302092 60088 302148
rect 269864 301420 279132 301476
rect 279188 301420 279198 301476
rect 55346 300860 55356 300916
rect 55412 300860 60116 300916
rect 54450 300748 54460 300804
rect 54516 300748 55356 300804
rect 55412 300748 55422 300804
rect 56690 300748 56700 300804
rect 56756 300748 57036 300804
rect 57092 300748 57102 300804
rect 60060 300776 60116 300860
rect 388098 300636 388108 300692
rect 388164 300636 476700 300692
rect 476756 300636 476766 300692
rect 388210 300524 388220 300580
rect 388276 300524 476476 300580
rect 476532 300524 476542 300580
rect 56914 300076 56924 300132
rect 56980 300076 60620 300132
rect 60676 300076 60686 300132
rect 269864 300076 277676 300132
rect 277732 300076 277742 300132
rect 56802 299404 56812 299460
rect 56868 299404 60088 299460
rect 269864 298732 270508 298788
rect 270564 298732 270574 298788
rect 57026 298060 57036 298116
rect 57092 298060 60088 298116
rect 595560 297892 597000 298088
rect 590818 297836 590828 297892
rect 590884 297864 597000 297892
rect 590884 297836 595672 297864
rect 269378 297388 269388 297444
rect 269444 297388 269454 297444
rect 388210 297276 388220 297332
rect 388276 297276 476812 297332
rect 476868 297276 476878 297332
rect 388434 297164 388444 297220
rect 388500 297164 476364 297220
rect 476420 297164 476430 297220
rect 60498 296716 60508 296772
rect 60564 296716 60574 296772
rect 56914 295372 56924 295428
rect 56980 295372 60088 295428
rect 56914 294028 56924 294084
rect 56980 294028 60088 294084
rect 476102 293916 476140 293972
rect 476196 293916 476206 293972
rect 56130 292684 56140 292740
rect 56196 292684 288316 292740
rect 288372 292684 288382 292740
rect 56466 292236 56476 292292
rect 56532 292236 293244 292292
rect 293300 292236 293310 292292
rect 388098 292236 388108 292292
rect 388164 292236 476252 292292
rect 476308 292236 476318 292292
rect 56578 292124 56588 292180
rect 56644 292124 289884 292180
rect 289940 292124 289950 292180
rect 56802 292012 56812 292068
rect 56868 292012 283052 292068
rect 283108 292012 283118 292068
rect 56354 291900 56364 291956
rect 56420 291900 281372 291956
rect 281428 291900 281438 291956
rect 56690 291788 56700 291844
rect 56756 291788 278236 291844
rect 278292 291788 278302 291844
rect 56242 291676 56252 291732
rect 56308 291676 276332 291732
rect 276388 291676 276398 291732
rect 56690 291564 56700 291620
rect 56756 291564 274652 291620
rect 274708 291564 274718 291620
rect 247762 291452 247772 291508
rect 247828 291452 272300 291508
rect 272356 291452 272366 291508
rect -960 290836 480 291032
rect -960 290808 4956 290836
rect 392 290780 4956 290808
rect 5012 290780 5022 290836
rect 388098 290556 388108 290612
rect 388164 290556 476588 290612
rect 476644 290556 476654 290612
rect 63718 290108 63756 290164
rect 63812 290108 63822 290164
rect 245186 289772 245196 289828
rect 245252 289772 269724 289828
rect 269780 289772 269790 289828
rect 475458 288988 475468 289044
rect 475524 288988 477036 289044
rect 477092 288988 477102 289044
rect 58146 288092 58156 288148
rect 58212 288092 115388 288148
rect 115444 288092 115454 288148
rect 180562 286972 180572 287028
rect 180628 286972 200284 287028
rect 200340 286972 200350 287028
rect 61170 286860 61180 286916
rect 61236 286860 103516 286916
rect 103572 286860 103582 286916
rect 155362 286860 155372 286916
rect 155428 286860 170044 286916
rect 170100 286860 170110 286916
rect 177202 286860 177212 286916
rect 177268 286860 210364 286916
rect 210420 286860 210430 286916
rect 26002 286748 26012 286804
rect 26068 286748 71260 286804
rect 71316 286748 71326 286804
rect 167122 286748 167132 286804
rect 167188 286748 206332 286804
rect 206388 286748 206398 286804
rect 27682 286636 27692 286692
rect 27748 286636 73276 286692
rect 73332 286636 73342 286692
rect 152002 286636 152012 286692
rect 152068 286636 194236 286692
rect 194292 286636 194302 286692
rect 58706 286524 58716 286580
rect 58772 286524 119644 286580
rect 119700 286524 119710 286580
rect 121762 286524 121772 286580
rect 121828 286524 131740 286580
rect 131796 286524 131806 286580
rect 143826 286524 143836 286580
rect 143892 286524 149660 286580
rect 149716 286524 149726 286580
rect 168802 286524 168812 286580
rect 168868 286524 212380 286580
rect 212436 286524 212446 286580
rect 59714 286412 59724 286468
rect 59780 286412 123676 286468
rect 123732 286412 123742 286468
rect 140242 286412 140252 286468
rect 140308 286412 190204 286468
rect 190260 286412 190270 286468
rect 200722 286412 200732 286468
rect 200788 286412 220444 286468
rect 220500 286412 220510 286468
rect 230962 286412 230972 286468
rect 231028 286412 236572 286468
rect 236628 286412 236638 286468
rect 254706 286412 254716 286468
rect 254772 286412 258748 286468
rect 258804 286412 258814 286468
rect 123442 286300 123452 286356
rect 123508 286300 127708 286356
rect 127764 286300 127774 286356
rect 135762 286300 135772 286356
rect 135828 286300 147980 286356
rect 148036 286300 148046 286356
rect 250674 286300 250684 286356
rect 250740 286300 255724 286356
rect 255780 286300 255790 286356
rect 136882 286188 136892 286244
rect 136948 286188 137788 286244
rect 137844 286188 137854 286244
rect 147858 286188 147868 286244
rect 147924 286188 149548 286244
rect 149604 286188 149614 286244
rect 145842 285964 145852 286020
rect 145908 285964 149772 286020
rect 149828 285964 149838 286020
rect 257954 285852 257964 285908
rect 258020 285852 262780 285908
rect 262836 285852 262846 285908
rect 149874 285740 149884 285796
rect 149940 285740 152908 285796
rect 152964 285740 152974 285796
rect 197362 285740 197372 285796
rect 197428 285740 202300 285796
rect 202356 285740 202366 285796
rect 227602 285740 227612 285796
rect 227668 285740 230524 285796
rect 230580 285740 230590 285796
rect 244626 285740 244636 285796
rect 244692 285740 252028 285796
rect 252084 285740 252094 285796
rect 259522 285740 259532 285796
rect 259588 285740 264796 285796
rect 264852 285740 264862 285796
rect 96562 285628 96572 285684
rect 96628 285628 97468 285684
rect 97524 285628 97534 285684
rect 124338 285628 124348 285684
rect 124404 285628 125692 285684
rect 125748 285628 125758 285684
rect 138562 285628 138572 285684
rect 138628 285628 139804 285684
rect 139860 285628 139870 285684
rect 141810 285628 141820 285684
rect 141876 285628 147868 285684
rect 147924 285628 147934 285684
rect 153010 285628 153020 285684
rect 153076 285628 153916 285684
rect 153972 285628 153982 285684
rect 154578 285628 154588 285684
rect 154644 285628 155932 285684
rect 155988 285628 155998 285684
rect 157042 285628 157052 285684
rect 157108 285628 157948 285684
rect 158004 285628 158014 285684
rect 159702 285628 159740 285684
rect 159796 285628 159806 285684
rect 164658 285628 164668 285684
rect 164724 285628 166012 285684
rect 166068 285628 166078 285684
rect 173058 285628 173068 285684
rect 173124 285628 174076 285684
rect 174132 285628 174142 285684
rect 174738 285628 174748 285684
rect 174804 285628 176092 285684
rect 176148 285628 176158 285684
rect 178070 285628 178108 285684
rect 178164 285628 178174 285684
rect 183138 285628 183148 285684
rect 183204 285628 184156 285684
rect 184212 285628 184222 285684
rect 184818 285628 184828 285684
rect 184884 285628 186172 285684
rect 186228 285628 186238 285684
rect 188150 285628 188188 285684
rect 188244 285628 188254 285684
rect 191510 285628 191548 285684
rect 191604 285628 191614 285684
rect 194898 285628 194908 285684
rect 194964 285628 196252 285684
rect 196308 285628 196318 285684
rect 198230 285628 198268 285684
rect 198324 285628 198334 285684
rect 203298 285628 203308 285684
rect 203364 285628 204316 285684
rect 204372 285628 204382 285684
rect 208338 285628 208348 285684
rect 208404 285628 208442 285684
rect 213378 285628 213388 285684
rect 213444 285628 214396 285684
rect 214452 285628 214462 285684
rect 215058 285628 215068 285684
rect 215124 285628 216412 285684
rect 216468 285628 216478 285684
rect 218390 285628 218428 285684
rect 218484 285628 218494 285684
rect 221750 285628 221788 285684
rect 221844 285628 221854 285684
rect 225138 285628 225148 285684
rect 225204 285628 226492 285684
rect 226548 285628 226558 285684
rect 228470 285628 228508 285684
rect 228564 285628 228574 285684
rect 231858 285628 231868 285684
rect 231924 285628 231962 285684
rect 237682 285628 237692 285684
rect 237748 285628 238588 285684
rect 238644 285628 238654 285684
rect 239362 285628 239372 285684
rect 239428 285628 240604 285684
rect 240660 285628 240670 285684
rect 242610 285628 242620 285684
rect 242676 285628 243516 285684
rect 243572 285628 243582 285684
rect 246838 285628 246876 285684
rect 246932 285628 246942 285684
rect 249190 285628 249228 285684
rect 249284 285628 249294 285684
rect 252102 285628 252140 285684
rect 252196 285628 252206 285684
rect 255602 285628 255612 285684
rect 255668 285628 256732 285684
rect 256788 285628 256798 285684
rect 257842 285628 257852 285684
rect 257908 285628 258748 285684
rect 258804 285628 258814 285684
rect 260390 285628 260428 285684
rect 260484 285628 260494 285684
rect 265458 285628 265468 285684
rect 265524 285628 266812 285684
rect 266868 285628 266878 285684
rect 29362 285068 29372 285124
rect 29428 285068 67228 285124
rect 67284 285068 67294 285124
rect 104962 285068 104972 285124
rect 105028 285068 151900 285124
rect 151956 285068 151966 285124
rect 49970 284956 49980 285012
rect 50036 284956 107324 285012
rect 107380 284956 107390 285012
rect 196018 284956 196028 285012
rect 196084 284956 270844 285012
rect 270900 284956 270910 285012
rect 58258 284844 58268 284900
rect 58324 284844 119420 284900
rect 119476 284844 119486 284900
rect 151666 284844 151676 284900
rect 151732 284844 270956 284900
rect 271012 284844 271022 284900
rect 590146 284844 590156 284900
rect 590212 284872 595672 284900
rect 590212 284844 597000 284872
rect 60162 284732 60172 284788
rect 60228 284732 135548 284788
rect 135604 284732 135614 284788
rect 143602 284732 143612 284788
rect 143668 284732 274092 284788
rect 274148 284732 274158 284788
rect 595560 284648 597000 284844
rect 51762 283276 51772 283332
rect 51828 283276 91196 283332
rect 91252 283276 91262 283332
rect 116722 283276 116732 283332
rect 116788 283276 163996 283332
rect 164052 283276 164062 283332
rect 200050 283276 200060 283332
rect 200116 283276 270732 283332
rect 270788 283276 270798 283332
rect 60274 283164 60284 283220
rect 60340 283164 127484 283220
rect 127540 283164 127550 283220
rect 191986 283164 191996 283220
rect 192052 283164 273980 283220
rect 274036 283164 274046 283220
rect 60050 283052 60060 283108
rect 60116 283052 139580 283108
rect 139636 283052 139646 283108
rect 147634 283052 147644 283108
rect 147700 283052 275660 283108
rect 275716 283052 275726 283108
rect 81442 281372 81452 281428
rect 81508 281372 115612 281428
rect 115668 281372 115678 281428
rect 171266 281372 171276 281428
rect 171332 281372 224476 281428
rect 224532 281372 224542 281428
rect 54898 281036 54908 281092
rect 54964 281036 476252 281092
rect 476308 281036 476318 281092
rect 54674 280700 54684 280756
rect 54740 280700 476476 280756
rect 476532 280700 476542 280756
rect 83122 280476 83132 280532
rect 83188 280476 473116 280532
rect 473172 280476 473182 280532
rect 83346 280364 83356 280420
rect 83412 280364 472892 280420
rect 472948 280364 472958 280420
rect 273746 279916 273756 279972
rect 273812 279916 304892 279972
rect 304948 279916 304958 279972
rect 273522 279804 273532 279860
rect 273588 279804 347788 279860
rect 347844 279804 347854 279860
rect 273074 279692 273084 279748
rect 273140 279692 355292 279748
rect 355348 279692 355358 279748
rect 374098 278796 374108 278852
rect 374164 278796 374444 278852
rect 374500 278796 374510 278852
rect 32722 278348 32732 278404
rect 32788 278348 81340 278404
rect 81396 278348 81406 278404
rect 273410 278348 273420 278404
rect 273476 278348 347900 278404
rect 347956 278348 347966 278404
rect 60610 278236 60620 278292
rect 60676 278236 565292 278292
rect 565348 278236 565358 278292
rect 60386 278124 60396 278180
rect 60452 278124 590604 278180
rect 590660 278124 590670 278180
rect 58258 278012 58268 278068
rect 58324 278012 590828 278068
rect 590884 278012 590894 278068
rect -960 276724 480 276920
rect 350242 276780 350252 276836
rect 350308 276780 375452 276836
rect 375508 276780 375518 276836
rect -960 276696 456092 276724
rect 392 276668 456092 276696
rect 456148 276668 456158 276724
rect 273186 276556 273196 276612
rect 273252 276556 350476 276612
rect 350532 276556 350542 276612
rect 56802 276444 56812 276500
rect 56868 276444 570332 276500
rect 570388 276444 570398 276500
rect 330866 276332 330876 276388
rect 330932 276332 419356 276388
rect 419412 276332 419422 276388
rect 308242 275660 308252 275716
rect 308308 275660 315868 275716
rect 315924 275660 315934 275716
rect 380482 275660 380492 275716
rect 380548 275660 384412 275716
rect 384468 275660 384478 275716
rect 309922 275548 309932 275604
rect 309988 275548 313292 275604
rect 313348 275548 313358 275604
rect 329634 275548 329644 275604
rect 329700 275548 330876 275604
rect 330932 275548 330942 275604
rect 352034 275548 352044 275604
rect 352100 275548 353948 275604
rect 354004 275548 354014 275604
rect 363794 275548 363804 275604
rect 363860 275548 366268 275604
rect 366324 275548 366334 275604
rect 382162 275548 382172 275604
rect 382228 275548 383516 275604
rect 383572 275548 383582 275604
rect 383842 275548 383852 275604
rect 383908 275548 385196 275604
rect 385252 275548 385262 275604
rect 273298 273196 273308 273252
rect 273364 273196 348012 273252
rect 348068 273196 348078 273252
rect 363122 273196 363132 273252
rect 363188 273196 385308 273252
rect 385364 273196 385374 273252
rect 56242 273084 56252 273140
rect 56308 273084 101500 273140
rect 101556 273084 101566 273140
rect 296482 273084 296492 273140
rect 296548 273084 580636 273140
rect 580692 273084 580702 273140
rect 58370 272972 58380 273028
rect 58436 272972 590492 273028
rect 590548 272972 590558 273028
rect 299842 271628 299852 271684
rect 299908 271628 454972 271684
rect 455028 271628 455038 271684
rect 4274 271516 4284 271572
rect 4340 271516 479612 271572
rect 479668 271516 479678 271572
rect 595560 271460 597000 271656
rect 74722 271404 74732 271460
rect 74788 271432 597000 271460
rect 74788 271404 595672 271432
rect 56914 271292 56924 271348
rect 56980 271292 566972 271348
rect 567028 271292 567038 271348
rect 248434 269948 248444 270004
rect 248500 269948 304444 270004
rect 304500 269948 304510 270004
rect 359426 269948 359436 270004
rect 359492 269948 390572 270004
rect 390628 269948 390638 270004
rect 56914 269836 56924 269892
rect 56980 269836 353612 269892
rect 353668 269836 353678 269892
rect 353938 269836 353948 269892
rect 354004 269836 396844 269892
rect 396900 269836 396910 269892
rect 4162 269724 4172 269780
rect 4228 269724 479612 269780
rect 479668 269724 479678 269780
rect 57026 269612 57036 269668
rect 57092 269612 568652 269668
rect 568708 269612 568718 269668
rect 356738 268268 356748 268324
rect 356804 268268 392812 268324
rect 392868 268268 392878 268324
rect 264562 268156 264572 268212
rect 264628 268156 364588 268212
rect 364644 268156 364654 268212
rect 366258 268156 366268 268212
rect 366324 268156 385084 268212
rect 385140 268156 385150 268212
rect 288194 268044 288204 268100
rect 288260 268044 590716 268100
rect 590772 268044 590782 268100
rect 56018 267932 56028 267988
rect 56084 267932 572012 267988
rect 572068 267932 572078 267988
rect 364466 266700 364476 266756
rect 364532 266700 380492 266756
rect 380548 266700 380558 266756
rect 356066 266588 356076 266644
rect 356132 266588 393372 266644
rect 393428 266588 393438 266644
rect 268594 266476 268604 266532
rect 268660 266476 371308 266532
rect 371364 266476 371374 266532
rect 50082 266364 50092 266420
rect 50148 266364 103292 266420
rect 103348 266364 103358 266420
rect 167794 266364 167804 266420
rect 167860 266364 269500 266420
rect 269556 266364 269566 266420
rect 289762 266364 289772 266420
rect 289828 266364 582540 266420
rect 582596 266364 582606 266420
rect 4498 266252 4508 266308
rect 4564 266252 477932 266308
rect 477988 266252 477998 266308
rect 363794 265132 363804 265188
rect 363860 265132 383852 265188
rect 383908 265132 383918 265188
rect 357746 265020 357756 265076
rect 357812 265020 391916 265076
rect 391972 265020 391982 265076
rect 276658 264908 276668 264964
rect 276724 264908 382172 264964
rect 382228 264908 382238 264964
rect 294914 264796 294924 264852
rect 294980 264796 584444 264852
rect 584500 264796 584510 264852
rect 4386 264684 4396 264740
rect 4452 264684 477932 264740
rect 477988 264684 477998 264740
rect 76402 264572 76412 264628
rect 76468 264572 590492 264628
rect 590548 264572 590558 264628
rect 374546 263004 374556 263060
rect 374612 263004 375452 263060
rect 375508 263004 375518 263060
rect 332434 262892 332444 262948
rect 332500 262892 417452 262948
rect 417508 262892 417518 262948
rect -960 262612 480 262808
rect 357074 262780 357084 262836
rect 357140 262780 365372 262836
rect 365428 262780 365438 262836
rect 373762 262780 373772 262836
rect 373828 262780 374556 262836
rect 374612 262780 374622 262836
rect 330306 262668 330316 262724
rect 330372 262668 418124 262724
rect 418180 262668 418190 262724
rect -960 262584 388892 262612
rect 392 262556 388892 262584
rect 388948 262556 388958 262612
rect 360322 262444 360332 262500
rect 360388 262444 373436 262500
rect 373492 262444 373502 262500
rect 374322 262444 374332 262500
rect 374388 262444 375004 262500
rect 375060 262444 375070 262500
rect 337652 262332 416332 262388
rect 416388 262332 416398 262388
rect 337652 262164 337708 262332
rect 374210 262220 374220 262276
rect 374276 262220 374668 262276
rect 374724 262220 374734 262276
rect 331762 262108 331772 262164
rect 331828 262108 332556 262164
rect 332612 262108 337708 262164
rect 372932 262108 376124 262164
rect 376180 262108 376190 262164
rect 372932 261492 372988 262108
rect 236338 261436 236348 261492
rect 236404 261436 372988 261492
rect 228274 261324 228284 261380
rect 228340 261324 423948 261380
rect 424004 261324 424014 261380
rect 55346 261212 55356 261268
rect 55412 261212 590716 261268
rect 590772 261212 590782 261268
rect 222562 260428 222572 260484
rect 222628 260428 435708 260484
rect 435764 260428 435774 260484
rect 224242 259756 224252 259812
rect 224308 259756 432236 259812
rect 432292 259756 432302 259812
rect 216178 259644 216188 259700
rect 216244 259644 443436 259700
rect 443492 259644 443502 259700
rect 73042 259532 73052 259588
rect 73108 259532 590604 259588
rect 590660 259532 590670 259588
rect 364214 259084 364252 259140
rect 364308 259084 364318 259140
rect 374966 259084 375004 259140
rect 375060 259084 375070 259140
rect 385718 259084 385756 259140
rect 385812 259084 385822 259140
rect 390534 259084 390572 259140
rect 390628 259084 390638 259140
rect 393894 259084 393932 259140
rect 393988 259084 393998 259140
rect 397254 259084 397292 259140
rect 397348 259084 397358 259140
rect 373846 258972 373884 259028
rect 373940 258972 373950 259028
rect 392214 258972 392252 259028
rect 392308 258972 392318 259028
rect 392438 258972 392476 259028
rect 392532 258972 392542 259028
rect 232306 258860 232316 258916
rect 232372 258860 384300 258916
rect 384356 258860 384366 258916
rect 385382 258860 385420 258916
rect 385476 258860 385486 258916
rect 208114 258748 208124 258804
rect 208180 258748 406588 258804
rect 406644 258748 406654 258804
rect 412374 258748 412412 258804
rect 412468 258748 412478 258804
rect 414054 258748 414092 258804
rect 414148 258748 414158 258804
rect 424358 258748 424396 258804
rect 424452 258748 424462 258804
rect 363878 258636 363916 258692
rect 363972 258636 363982 258692
rect 373762 258636 373772 258692
rect 373828 258636 374332 258692
rect 374388 258636 374398 258692
rect 374882 258636 374892 258692
rect 374948 258636 375228 258692
rect 375284 258636 375294 258692
rect 433458 258636 433468 258692
rect 433524 258636 434924 258692
rect 434980 258636 434990 258692
rect 433794 258524 433804 258580
rect 433860 258524 434252 258580
rect 434308 258524 434318 258580
rect 423378 258412 423388 258468
rect 423444 258412 424060 258468
rect 424116 258412 424126 258468
rect 434102 258412 434140 258468
rect 434196 258412 434206 258468
rect 434550 258412 434588 258468
rect 434644 258412 434654 258468
rect 444630 258412 444668 258468
rect 444724 258412 444734 258468
rect 445302 258412 445340 258468
rect 445396 258412 445406 258468
rect 595560 258244 597000 258440
rect 572002 258188 572012 258244
rect 572068 258216 597000 258244
rect 572068 258188 595672 258216
rect 86482 257964 86492 258020
rect 86548 257964 129724 258020
rect 129780 257964 129790 258020
rect 48402 257852 48412 257908
rect 48468 257852 99260 257908
rect 99316 257852 99326 257908
rect 204082 257852 204092 257908
rect 204148 257852 270620 257908
rect 270676 257852 270686 257908
rect 272962 257852 272972 257908
rect 273028 257852 356972 257908
rect 357028 257852 357038 257908
rect 45602 254492 45612 254548
rect 45668 254492 93436 254548
rect 93492 254492 93502 254548
rect 240370 254492 240380 254548
rect 240436 254492 360332 254548
rect 360388 254492 360398 254548
rect 34402 252812 34412 252868
rect 34468 252812 83356 252868
rect 83412 252812 83422 252868
rect 42802 251132 42812 251188
rect 42868 251132 91420 251188
rect 91476 251132 91486 251188
rect -960 248500 480 248696
rect -960 248472 4172 248500
rect 392 248444 4172 248472
rect 4228 248444 4238 248500
rect 49522 246092 49532 246148
rect 49588 246092 95452 246148
rect 95508 246092 95518 246148
rect 590706 245196 590716 245252
rect 590772 245224 595672 245252
rect 590772 245196 597000 245224
rect 595560 245000 597000 245196
rect 392 234584 4172 234612
rect -960 234556 4172 234584
rect 4228 234556 4238 234612
rect -960 234360 480 234556
rect 51202 234332 51212 234388
rect 51268 234332 85372 234388
rect 85428 234332 85438 234388
rect 44482 232652 44492 232708
rect 44548 232652 89404 232708
rect 89460 232652 89470 232708
rect 590818 231980 590828 232036
rect 590884 232008 595672 232036
rect 590884 231980 597000 232008
rect 595560 231784 597000 231980
rect 89842 231084 89852 231140
rect 89908 231084 133756 231140
rect 133812 231084 133822 231140
rect 24322 230972 24332 231028
rect 24388 230972 69244 231028
rect 69300 230972 69310 231028
rect 133522 230972 133532 231028
rect 133588 230972 180124 231028
rect 180180 230972 180190 231028
rect 53218 229292 53228 229348
rect 53284 229292 99484 229348
rect 99540 229292 99550 229348
rect 70354 227724 70364 227780
rect 70420 227724 117628 227780
rect 117684 227724 117694 227780
rect 50194 227612 50204 227668
rect 50260 227612 123452 227668
rect 123508 227612 123518 227668
rect 37986 224252 37996 224308
rect 38052 224252 87388 224308
rect 87444 224252 87454 224308
rect 187954 224252 187964 224308
rect 188020 224252 275548 224308
rect 275604 224252 275614 224308
rect 48514 222684 48524 222740
rect 48580 222684 87164 222740
rect 87220 222684 87230 222740
rect 260530 222684 260540 222740
rect 260596 222684 322588 222740
rect 322644 222684 322654 222740
rect 49410 222572 49420 222628
rect 49476 222572 96572 222628
rect 96628 222572 96638 222628
rect 109106 222572 109116 222628
rect 109172 222572 157052 222628
rect 157108 222572 157118 222628
rect 163762 222572 163772 222628
rect 163828 222572 270508 222628
rect 270564 222572 270574 222628
rect 392 220472 4508 220500
rect -960 220444 4508 220472
rect 4564 220444 4574 220500
rect -960 220248 480 220444
rect 47842 219212 47852 219268
rect 47908 219212 79324 219268
rect 79380 219212 79390 219268
rect 590706 218764 590716 218820
rect 590772 218792 595672 218820
rect 590772 218764 597000 218792
rect 595560 218568 597000 218764
rect 24658 217644 24668 217700
rect 24724 217644 77308 217700
rect 77364 217644 77374 217700
rect 244402 217644 244412 217700
rect 244468 217644 357084 217700
rect 357140 217644 357150 217700
rect 58370 217532 58380 217588
rect 58436 217532 131516 217588
rect 131572 217532 131582 217588
rect 155698 217532 155708 217588
rect 155764 217532 269388 217588
rect 269444 217532 269454 217588
rect 256498 215964 256508 216020
rect 256564 215964 308252 216020
rect 308308 215964 308318 216020
rect 48626 215852 48636 215908
rect 48692 215852 111356 215908
rect 111412 215852 111422 215908
rect 212146 215852 212156 215908
rect 212212 215852 342636 215908
rect 342692 215852 342702 215908
rect 31042 214284 31052 214340
rect 31108 214284 75292 214340
rect 75348 214284 75358 214340
rect 252466 214284 252476 214340
rect 252532 214284 309932 214340
rect 309988 214284 309998 214340
rect 58594 214172 58604 214228
rect 58660 214172 121660 214228
rect 121716 214172 121726 214228
rect 183922 214172 183932 214228
rect 183988 214172 273868 214228
rect 273924 214172 273934 214228
rect 66630 213276 66668 213332
rect 66724 213276 66734 213332
rect 220210 213276 220220 213332
rect 220276 213276 222572 213332
rect 222628 213276 222638 213332
rect 59826 212940 59836 212996
rect 59892 212940 75068 212996
rect 75124 212940 75134 212996
rect 55234 212828 55244 212884
rect 55300 212828 71036 212884
rect 71092 212828 71102 212884
rect 179890 212828 179900 212884
rect 179956 212828 271516 212884
rect 271572 212828 271582 212884
rect 59602 212716 59612 212772
rect 59668 212716 83132 212772
rect 83188 212716 83198 212772
rect 130162 212716 130172 212772
rect 130228 212716 172060 212772
rect 172116 212716 172126 212772
rect 175858 212716 175868 212772
rect 175924 212716 269836 212772
rect 269892 212716 269902 212772
rect 53666 212604 53676 212660
rect 53732 212604 79100 212660
rect 79156 212604 79166 212660
rect 171826 212604 171836 212660
rect 171892 212604 271292 212660
rect 271348 212604 271358 212660
rect 60610 212492 60620 212548
rect 60676 212492 95228 212548
rect 95284 212492 95294 212548
rect 159730 212492 159740 212548
rect 159796 212492 269612 212548
rect 269668 212492 269678 212548
rect 272626 212492 272636 212548
rect 272692 212492 350252 212548
rect 350308 212492 350318 212548
rect 58930 211148 58940 211204
rect 58996 211148 105532 211204
rect 105588 211148 105598 211204
rect 17602 211036 17612 211092
rect 17668 211036 65212 211092
rect 65268 211036 65278 211092
rect 60274 210924 60284 210980
rect 60340 210924 111580 210980
rect 111636 210924 111646 210980
rect 135202 210924 135212 210980
rect 135268 210924 182140 210980
rect 182196 210924 182206 210980
rect 60162 210812 60172 210868
rect 60228 210812 113596 210868
rect 113652 210812 113662 210868
rect 119186 210812 119196 210868
rect 119252 210812 168028 210868
rect 168084 210812 168094 210868
rect 182242 210812 182252 210868
rect 182308 210812 234556 210868
rect 234612 210812 234622 210868
rect 62934 209916 62972 209972
rect 63028 209916 63038 209972
rect 59938 209468 59948 209524
rect 60004 209468 107548 209524
rect 107604 209468 107614 209524
rect 60050 209356 60060 209412
rect 60116 209356 109564 209412
rect 109620 209356 109630 209412
rect 112466 209356 112476 209412
rect 112532 209356 161980 209412
rect 162036 209356 162046 209412
rect 392 206360 4172 206388
rect -960 206332 4172 206360
rect 4228 206332 4238 206388
rect -960 206136 480 206332
rect 590146 205548 590156 205604
rect 590212 205576 595672 205604
rect 590212 205548 597000 205576
rect 595560 205352 597000 205548
rect 590594 192332 590604 192388
rect 590660 192360 595672 192388
rect 590660 192332 597000 192360
rect 392 192248 4396 192276
rect -960 192220 4396 192248
rect 4452 192220 4462 192276
rect -960 192024 480 192220
rect 595560 192136 597000 192332
rect 595560 178948 597000 179144
rect 570322 178892 570332 178948
rect 570388 178920 597000 178948
rect 570388 178892 595672 178920
rect -960 178052 480 178136
rect -960 177996 4284 178052
rect 4340 177996 4350 178052
rect -960 177912 480 177996
rect 284722 170492 284732 170548
rect 284788 170492 357868 170548
rect 357924 170492 357934 170548
rect 298162 168812 298172 168868
rect 298228 168812 352156 168868
rect 352212 168812 352222 168868
rect 590594 165900 590604 165956
rect 590660 165928 595672 165956
rect 590660 165900 597000 165928
rect 595560 165704 597000 165900
rect 392 164024 4172 164052
rect -960 163996 4172 164024
rect 4228 163996 4238 164052
rect -960 163800 480 163996
rect 293122 163772 293132 163828
rect 293188 163772 329308 163828
rect 329364 163772 329374 163828
rect 291442 162092 291452 162148
rect 291508 162092 322588 162148
rect 322644 162092 322654 162148
rect 4162 160636 4172 160692
rect 4228 160636 467852 160692
rect 467908 160636 467918 160692
rect 60498 160524 60508 160580
rect 60564 160524 590828 160580
rect 590884 160524 590894 160580
rect 51986 160412 51996 160468
rect 52052 160412 590604 160468
rect 590660 160412 590670 160468
rect 233426 160300 233436 160356
rect 233492 160300 279132 160356
rect 279188 160300 279198 160356
rect 267026 160188 267036 160244
rect 267092 160188 279020 160244
rect 279076 160188 279086 160244
rect 501218 160076 501228 160132
rect 501284 160076 502124 160132
rect 502180 160076 502190 160132
rect 483970 159628 483980 159684
rect 484036 159628 485212 159684
rect 485268 159628 485278 159684
rect 146962 159516 146972 159572
rect 147028 159516 512316 159572
rect 512372 159516 512382 159572
rect 257170 159404 257180 159460
rect 257236 159404 475020 159460
rect 475076 159404 475086 159460
rect 226706 158956 226716 159012
rect 226772 158956 277676 159012
rect 277732 158956 277742 159012
rect 468626 158956 468636 159012
rect 468692 158956 552076 159012
rect 552132 158956 552142 159012
rect 80546 158844 80556 158900
rect 80612 158844 123452 158900
rect 123508 158844 123518 158900
rect 157266 158844 157276 158900
rect 157332 158844 191548 158900
rect 191604 158844 191614 158900
rect 260418 158844 260428 158900
rect 260484 158844 267148 158900
rect 273858 158844 273868 158900
rect 273924 158844 485884 158900
rect 485940 158844 485950 158900
rect 267092 158788 267148 158844
rect 78866 158732 78876 158788
rect 78932 158732 124348 158788
rect 124404 158732 124414 158788
rect 179666 158732 179676 158788
rect 179732 158732 231868 158788
rect 231924 158732 231934 158788
rect 267092 158732 483196 158788
rect 483252 158732 483262 158788
rect 262546 157836 262556 157892
rect 262612 157836 273868 157892
rect 273924 157836 273934 157892
rect 275986 157836 275996 157892
rect 276052 157836 553532 157892
rect 553588 157836 553598 157892
rect 69010 157724 69020 157780
rect 69076 157724 73836 157780
rect 73892 157724 73902 157780
rect 270610 157724 270620 157780
rect 270676 157724 542892 157780
rect 542948 157724 542958 157780
rect 273298 157612 273308 157668
rect 273364 157612 545468 157668
rect 545524 157612 545534 157668
rect 216850 157500 216860 157556
rect 216916 157500 252812 157556
rect 252868 157500 252878 157556
rect 265234 157500 265244 157556
rect 265300 157500 493948 157556
rect 494004 157500 494014 157556
rect 208786 157388 208796 157444
rect 208852 157388 247772 157444
rect 247828 157388 247838 157444
rect 117394 157276 117404 157332
rect 117460 157276 133756 157332
rect 133812 157276 133822 157332
rect 149090 157276 149100 157332
rect 149156 157276 160412 157332
rect 160468 157276 160478 157332
rect 179218 157276 179228 157332
rect 179284 157276 222572 157332
rect 222628 157276 222638 157332
rect 254482 157276 254492 157332
rect 254548 157276 265468 157332
rect 265524 157276 265534 157332
rect 74386 157164 74396 157220
rect 74452 157164 123564 157220
rect 123620 157164 123630 157220
rect 146962 157164 146972 157220
rect 147028 157164 165788 157220
rect 165844 157164 165854 157220
rect 195346 157164 195356 157220
rect 195412 157164 241948 157220
rect 242004 157164 242014 157220
rect 246418 157164 246428 157220
rect 246484 157164 261212 157220
rect 261268 157164 261278 157220
rect 71698 157052 71708 157108
rect 71764 157052 133980 157108
rect 134036 157052 134046 157108
rect 155362 157052 155372 157108
rect 155428 157052 184828 157108
rect 184884 157052 184894 157108
rect 192658 157052 192668 157108
rect 192724 157052 246652 157108
rect 246708 157052 246718 157108
rect 249106 157052 249116 157108
rect 249172 157052 264572 157108
rect 264628 157052 264638 157108
rect 267922 157052 267932 157108
rect 267988 157052 308252 157108
rect 308308 157052 308318 157108
rect 66322 156492 66332 156548
rect 66388 156492 70476 156548
rect 70532 156492 70542 156548
rect 230290 156492 230300 156548
rect 230356 156492 234332 156548
rect 234388 156492 234398 156548
rect 153682 156268 153692 156324
rect 153748 156268 155036 156324
rect 155092 156268 155102 156324
rect 162082 156268 162092 156324
rect 162148 156268 163100 156324
rect 163156 156268 163166 156324
rect 188962 156268 188972 156324
rect 189028 156268 189980 156324
rect 190036 156268 190046 156324
rect 243730 156268 243740 156324
rect 243796 156268 246092 156324
rect 246148 156268 246158 156324
rect 251794 156268 251804 156324
rect 251860 156268 258636 156324
rect 258692 156268 258702 156324
rect 474534 156268 474572 156324
rect 474628 156268 474638 156324
rect 308242 156156 308252 156212
rect 308308 156156 534604 156212
rect 534660 156156 534670 156212
rect 200722 155820 200732 155876
rect 200788 155820 324940 155876
rect 324996 155820 325006 155876
rect 93202 155708 93212 155764
rect 93268 155708 116732 155764
rect 116788 155708 116798 155764
rect 138898 155708 138908 155764
rect 138964 155708 306572 155764
rect 306628 155708 306638 155764
rect 106642 155596 106652 155652
rect 106708 155596 133532 155652
rect 133588 155596 133598 155652
rect 258626 155596 258636 155652
rect 258692 155596 473452 155652
rect 473508 155596 473518 155652
rect 493042 155596 493052 155652
rect 493108 155596 526092 155652
rect 526148 155596 526158 155652
rect 63858 155484 63868 155540
rect 63924 155484 96908 155540
rect 96964 155484 96974 155540
rect 112018 155484 112028 155540
rect 112084 155484 144508 155540
rect 144564 155484 144574 155540
rect 214162 155484 214172 155540
rect 214228 155484 443884 155540
rect 443940 155484 443950 155540
rect 491362 155484 491372 155540
rect 491428 155484 527996 155540
rect 528052 155484 528062 155540
rect 73826 155372 73836 155428
rect 73892 155372 134652 155428
rect 134708 155372 134718 155428
rect 141586 155372 141596 155428
rect 141652 155372 406588 155428
rect 406644 155372 406654 155428
rect 464706 155372 464716 155428
rect 464772 155372 555100 155428
rect 555156 155372 555166 155428
rect 225138 153692 225148 153748
rect 225204 153692 384412 153748
rect 384468 153692 384478 153748
rect 176082 152796 176092 152852
rect 176148 152796 184604 152852
rect 184660 152796 184670 152852
rect 595560 152516 597000 152712
rect 58034 152460 58044 152516
rect 58100 152488 597000 152516
rect 58100 152460 595672 152488
rect 160850 152348 160860 152404
rect 160916 152348 228508 152404
rect 228564 152348 228574 152404
rect 255042 152348 255052 152404
rect 255108 152348 278908 152404
rect 278964 152348 278974 152404
rect 203410 152236 203420 152292
rect 203476 152236 284284 152292
rect 284340 152236 284350 152292
rect 294802 152236 294812 152292
rect 294868 152236 449260 152292
rect 449316 152236 449326 152292
rect 486322 152236 486332 152292
rect 486388 152236 533148 152292
rect 533204 152236 533214 152292
rect 70466 152124 70476 152180
rect 70532 152124 144732 152180
rect 144788 152124 144798 152180
rect 222226 152124 222236 152180
rect 222292 152124 424956 152180
rect 425012 152124 425022 152180
rect 474562 152124 474572 152180
rect 474628 152124 544348 152180
rect 544404 152124 544414 152180
rect 144274 152012 144284 152068
rect 144340 152012 506604 152068
rect 506660 152012 506670 152068
rect 257842 151116 257852 151172
rect 257908 151116 265468 151172
rect 265524 151116 265534 151172
rect 241938 150668 241948 150724
rect 242004 150668 335692 150724
rect 335748 150668 335758 150724
rect 155474 150556 155484 150612
rect 155540 150556 188188 150612
rect 188244 150556 188254 150612
rect 198258 150556 198268 150612
rect 198324 150556 333116 150612
rect 333172 150556 333182 150612
rect 491586 150556 491596 150612
rect 491652 150556 526988 150612
rect 527044 150556 527054 150612
rect 174738 150444 174748 150500
rect 174804 150444 235788 150500
rect 235844 150444 235854 150500
rect 265458 150444 265468 150500
rect 265524 150444 465388 150500
rect 465444 150444 465454 150500
rect 475458 150444 475468 150500
rect 475524 150444 542556 150500
rect 542612 150444 542622 150500
rect 65426 150332 65436 150388
rect 65492 150332 168476 150388
rect 168532 150332 168542 150388
rect 219538 150332 219548 150388
rect 219604 150332 433132 150388
rect 433188 150332 433198 150388
rect 464482 150332 464492 150388
rect 464548 150332 554316 150388
rect 554372 150332 554382 150388
rect -960 149716 480 149912
rect -960 149688 462812 149716
rect 392 149660 462812 149688
rect 462868 149660 462878 149716
rect 260306 148764 260316 148820
rect 260372 148764 272188 148820
rect 272244 148764 272254 148820
rect 77074 148652 77084 148708
rect 77140 148652 85036 148708
rect 85092 148652 85102 148708
rect 109330 148652 109340 148708
rect 109396 148652 118188 148708
rect 118244 148652 118254 148708
rect 148418 148652 148428 148708
rect 148484 148652 180572 148708
rect 180628 148652 180638 148708
rect 249330 148652 249340 148708
rect 249396 148652 278796 148708
rect 278852 148652 278862 148708
rect 120082 147868 120092 147924
rect 120148 147868 123340 147924
rect 123396 147868 123406 147924
rect 181906 147868 181916 147924
rect 181972 147868 184268 147924
rect 184324 147868 184334 147924
rect 247762 147420 247772 147476
rect 247828 147420 273420 147476
rect 273476 147420 273486 147476
rect 211474 147308 211484 147364
rect 211540 147308 265356 147364
rect 265412 147308 265422 147364
rect 150322 147196 150332 147252
rect 150388 147196 197372 147252
rect 197428 147196 197438 147252
rect 246642 147196 246652 147252
rect 246708 147196 343868 147252
rect 343924 147196 343934 147252
rect 106754 147084 106764 147140
rect 106820 147084 117516 147140
rect 117572 147084 117582 147140
rect 157490 147084 157500 147140
rect 157556 147084 164668 147140
rect 164724 147084 164734 147140
rect 176530 147084 176540 147140
rect 176596 147084 233100 147140
rect 233156 147084 233166 147140
rect 252802 147084 252812 147140
rect 252868 147084 435708 147140
rect 435764 147084 435774 147140
rect 474114 147084 474124 147140
rect 474180 147084 544572 147140
rect 544628 147084 544638 147140
rect 76066 146972 76076 147028
rect 76132 146972 162092 147028
rect 162148 146972 162158 147028
rect 171154 146972 171164 147028
rect 171220 146972 243852 147028
rect 243908 146972 243918 147028
rect 264562 146972 264572 147028
rect 264628 146972 476028 147028
rect 476084 146972 476094 147028
rect 493378 146972 493388 147028
rect 493444 146972 524188 147028
rect 524244 146972 524254 147028
rect 246866 146188 246876 146244
rect 246932 146188 247548 146244
rect 247604 146188 247614 146244
rect 150434 145740 150444 145796
rect 150500 145740 174748 145796
rect 174804 145740 174814 145796
rect 232978 145740 232988 145796
rect 233044 145740 365372 145796
rect 365428 145740 365438 145796
rect 496850 145740 496860 145796
rect 496916 145740 520828 145796
rect 520884 145740 520894 145796
rect 125010 145628 125020 145684
rect 125076 145628 157724 145684
rect 157780 145628 157790 145684
rect 159842 145628 159852 145684
rect 159908 145628 168812 145684
rect 168868 145628 168878 145684
rect 173506 145628 173516 145684
rect 173572 145628 187292 145684
rect 187348 145628 187358 145684
rect 227602 145628 227612 145684
rect 227668 145628 376124 145684
rect 376180 145628 376190 145684
rect 475010 145628 475020 145684
rect 475076 145628 542668 145684
rect 542724 145628 542734 145684
rect 90514 145516 90524 145572
rect 90580 145516 114716 145572
rect 114772 145516 114782 145572
rect 136210 145516 136220 145572
rect 136276 145516 206556 145572
rect 206612 145516 206622 145572
rect 241042 145516 241052 145572
rect 241108 145516 533036 145572
rect 533092 145516 533102 145572
rect 73490 145404 73500 145460
rect 73556 145404 146972 145460
rect 147028 145404 147038 145460
rect 152002 145404 152012 145460
rect 152068 145404 194908 145460
rect 194964 145404 194974 145460
rect 238354 145404 238364 145460
rect 238420 145404 535724 145460
rect 535780 145404 535790 145460
rect 55234 145292 55244 145348
rect 55300 145292 590604 145348
rect 590660 145292 590670 145348
rect 143826 144396 143836 144452
rect 143892 144396 149660 144452
rect 149716 144396 149726 144452
rect 154130 144172 154140 144228
rect 154196 144172 167132 144228
rect 167188 144172 167198 144228
rect 133074 144060 133084 144116
rect 133140 144060 153692 144116
rect 153748 144060 153758 144116
rect 165330 144060 165340 144116
rect 165396 144060 188972 144116
rect 189028 144060 189038 144116
rect 206098 144060 206108 144116
rect 206164 144060 276108 144116
rect 276164 144060 276174 144116
rect 315410 144060 315420 144116
rect 315476 144060 315756 144116
rect 315812 144060 315822 144116
rect 148642 143948 148652 144004
rect 148708 143948 173068 144004
rect 173124 143948 173134 144004
rect 222562 143948 222572 144004
rect 222628 143948 224924 144004
rect 224980 143948 224990 144004
rect 234322 143948 234332 144004
rect 234388 143948 373436 144004
rect 373492 143948 373502 144004
rect 148866 143836 148876 143892
rect 148932 143836 178108 143892
rect 178164 143836 178174 143892
rect 243506 143836 243516 143892
rect 243572 143836 250348 143892
rect 250404 143836 250414 143892
rect 261202 143836 261212 143892
rect 261268 143836 484316 143892
rect 484372 143836 484382 143892
rect 485090 143836 485100 143892
rect 485156 143836 532588 143892
rect 532644 143836 532654 143892
rect 87826 143724 87836 143780
rect 87892 143724 112588 143780
rect 112644 143724 112654 143780
rect 114706 143724 114716 143780
rect 114772 143724 134988 143780
rect 135044 143724 135054 143780
rect 135650 143724 135660 143780
rect 135716 143724 152348 143780
rect 152404 143724 152414 143780
rect 152562 143724 152572 143780
rect 152628 143724 183148 143780
rect 183204 143724 183214 143780
rect 246082 143724 246092 143780
rect 246148 143724 524972 143780
rect 525028 143724 525038 143780
rect 84242 143612 84252 143668
rect 84308 143612 149100 143668
rect 149156 143612 149166 143668
rect 157938 143612 157948 143668
rect 158004 143612 177212 143668
rect 177268 143612 177278 143668
rect 180562 143612 180572 143668
rect 180628 143612 225148 143668
rect 225204 143612 225214 143668
rect 235666 143612 235676 143668
rect 235732 143612 543900 143668
rect 543956 143612 543966 143668
rect 315522 143276 315532 143332
rect 315588 143276 334124 143332
rect 334180 143276 334190 143332
rect 315410 143164 315420 143220
rect 315476 143164 333788 143220
rect 333844 143164 333854 143220
rect 315746 143052 315756 143108
rect 315812 143052 334572 143108
rect 334628 143052 334638 143108
rect 312498 142940 312508 142996
rect 312564 142940 314076 142996
rect 314132 142940 335020 142996
rect 335076 142940 335086 142996
rect 495394 142940 495404 142996
rect 495460 142940 523404 142996
rect 523460 142940 523470 142996
rect 314132 142828 334348 142884
rect 334404 142828 334414 142884
rect 498978 142828 498988 142884
rect 499044 142828 500556 142884
rect 500612 142828 519260 142884
rect 519316 142828 519326 142884
rect 144694 142716 144732 142772
rect 144788 142716 144798 142772
rect 304742 142716 304780 142772
rect 304836 142716 304846 142772
rect 129266 142604 129276 142660
rect 129332 142604 174188 142660
rect 174244 142604 174254 142660
rect 112578 142492 112588 142548
rect 112644 142492 196588 142548
rect 196532 142436 196588 142492
rect 314132 142436 314188 142828
rect 330838 142716 330876 142772
rect 330932 142716 330942 142772
rect 333414 142716 333452 142772
rect 333508 142716 333518 142772
rect 412374 142716 412412 142772
rect 412468 142716 412478 142772
rect 463810 142716 463820 142772
rect 463876 142716 464716 142772
rect 464772 142716 464782 142772
rect 385522 142604 385532 142660
rect 385588 142604 485100 142660
rect 485156 142604 485166 142660
rect 375106 142492 375116 142548
rect 375172 142492 475020 142548
rect 475076 142492 475086 142548
rect 144498 142380 144508 142436
rect 144564 142380 145404 142436
rect 145460 142380 145470 142436
rect 196532 142380 212940 142436
rect 212996 142380 312956 142436
rect 313012 142380 314188 142436
rect 323810 142380 323820 142436
rect 323876 142380 325052 142436
rect 325108 142380 423724 142436
rect 423780 142380 423790 142436
rect 433682 142380 433692 142436
rect 433748 142380 478828 142436
rect 64418 142268 64428 142324
rect 64484 142268 84924 142324
rect 84980 142268 84990 142324
rect 130918 142268 130956 142324
rect 131012 142268 163772 142324
rect 163828 142268 164556 142324
rect 164612 142268 164622 142324
rect 234994 142268 235004 142324
rect 235060 142268 315756 142324
rect 315812 142268 315822 142324
rect 316418 142268 316428 142324
rect 316484 142268 331772 142324
rect 331828 142268 331838 142324
rect 364214 142268 364252 142324
rect 364308 142268 364318 142324
rect 364466 142268 364476 142324
rect 364532 142268 464492 142324
rect 464548 142268 464558 142324
rect 74610 142156 74620 142212
rect 74676 142156 82460 142212
rect 82516 142156 174636 142212
rect 174692 142156 174702 142212
rect 235106 142156 235116 142212
rect 235172 142156 315532 142212
rect 315588 142156 315598 142212
rect 364252 142100 364308 142268
rect 374546 142156 374556 142212
rect 374612 142156 474572 142212
rect 474628 142156 474638 142212
rect 478772 142100 478828 142380
rect 498978 142268 498988 142324
rect 499044 142268 501452 142324
rect 501508 142268 517468 142324
rect 517524 142268 517534 142324
rect 495506 142156 495516 142212
rect 495572 142156 523740 142212
rect 523796 142156 523806 142212
rect 75058 142044 75068 142100
rect 75124 142044 79772 142100
rect 79828 142044 174972 142100
rect 175028 142044 176316 142100
rect 176372 142044 176382 142100
rect 186386 142044 186396 142100
rect 186452 142044 285068 142100
rect 285124 142044 285134 142100
rect 317426 142044 317436 142100
rect 317492 142044 332444 142100
rect 332500 142044 336028 142100
rect 336084 142044 336094 142100
rect 344614 142044 344652 142100
rect 344708 142044 344718 142100
rect 364252 142044 463820 142100
rect 463876 142044 463886 142100
rect 478772 142044 484652 142100
rect 484708 142044 534156 142100
rect 534212 142044 534222 142100
rect 11330 141932 11340 141988
rect 11396 141932 62188 141988
rect 62244 141932 62254 141988
rect 74162 141932 74172 141988
rect 74228 141932 128156 141988
rect 128212 141932 129276 141988
rect 129332 141932 129342 141988
rect 164546 141932 164556 141988
rect 164612 141932 263788 141988
rect 263844 141932 263854 141988
rect 334114 141932 334124 141988
rect 334180 141932 433692 141988
rect 433748 141932 434140 141988
rect 434196 141932 434206 141988
rect 444630 141932 444668 141988
rect 444724 141932 444734 141988
rect 471986 141932 471996 141988
rect 472052 141932 472892 141988
rect 472948 141932 545356 141988
rect 545412 141932 545422 141988
rect 134642 141820 134652 141876
rect 134708 141820 234556 141876
rect 234612 141820 235004 141876
rect 235060 141820 235070 141876
rect 264450 141820 264460 141876
rect 264516 141820 363692 141876
rect 363748 141820 364476 141876
rect 364532 141820 364542 141876
rect 373314 141820 373324 141876
rect 373380 141820 375004 141876
rect 375060 141820 375116 141876
rect 375172 141820 375182 141876
rect 423714 141820 423724 141876
rect 423780 141820 424396 141876
rect 424452 141820 494732 141876
rect 494788 141820 495516 141876
rect 495572 141820 495582 141876
rect 90962 141708 90972 141764
rect 91028 141708 95900 141764
rect 95956 141708 96460 141764
rect 96516 141708 96526 141764
rect 176306 141708 176316 141764
rect 176372 141708 274988 141764
rect 275044 141708 275054 141764
rect 318210 141708 318220 141764
rect 318276 141708 330316 141764
rect 330372 141708 330876 141764
rect 330932 141708 330942 141764
rect 334338 141708 334348 141764
rect 334404 141708 412412 141764
rect 412468 141708 420028 141764
rect 433794 141708 433804 141764
rect 433860 141708 434364 141764
rect 434420 141708 434430 141764
rect 434578 141708 434588 141764
rect 434644 141708 484092 141764
rect 484148 141708 484428 141764
rect 484484 141708 484494 141764
rect 484866 141708 484876 141764
rect 484932 141708 485436 141764
rect 485492 141708 534940 141764
rect 534996 141708 535006 141764
rect 419972 141652 420028 141708
rect 174626 141596 174636 141652
rect 174692 141596 274540 141652
rect 274596 141596 373436 141652
rect 373492 141596 373502 141652
rect 373660 141596 384748 141652
rect 419972 141596 507276 141652
rect 507332 141596 512988 141652
rect 513044 141596 513054 141652
rect 373660 141540 373716 141596
rect 91970 141484 91980 141540
rect 92036 141484 97692 141540
rect 97748 141484 98588 141540
rect 98644 141484 98654 141540
rect 123554 141484 123564 141540
rect 123620 141484 223804 141540
rect 223860 141484 323820 141540
rect 323876 141484 323886 141540
rect 334562 141484 334572 141540
rect 334628 141484 373716 141540
rect 384692 141540 384748 141596
rect 384692 141484 434588 141540
rect 434644 141484 434654 141540
rect 505558 141484 505596 141540
rect 505652 141484 514668 141540
rect 514724 141484 514734 141540
rect 85810 141372 85820 141428
rect 85876 141372 122668 141428
rect 122724 141372 122734 141428
rect 133970 141372 133980 141428
rect 134036 141372 234220 141428
rect 234276 141372 235116 141428
rect 235172 141372 235182 141428
rect 274978 141372 274988 141428
rect 275044 141372 373324 141428
rect 373380 141372 373390 141428
rect 374770 141372 374780 141428
rect 374836 141372 375452 141428
rect 375508 141372 375518 141428
rect 503906 141372 503916 141428
rect 503972 141372 516348 141428
rect 516404 141372 516414 141428
rect 75506 141260 75516 141316
rect 75572 141260 124348 141316
rect 124404 141260 124414 141316
rect 164406 141260 164444 141316
rect 164500 141260 264460 141316
rect 264516 141260 264526 141316
rect 285058 141260 285068 141316
rect 285124 141260 385084 141316
rect 385140 141260 385532 141316
rect 385588 141260 385598 141316
rect 500658 141260 500668 141316
rect 500724 141260 502236 141316
rect 502292 141260 518140 141316
rect 518196 141260 518206 141316
rect 63718 141148 63756 141204
rect 63812 141148 63822 141204
rect 92754 141148 92764 141204
rect 92820 141148 100828 141204
rect 100884 141148 100894 141204
rect 114678 141148 114716 141204
rect 114772 141148 114782 141204
rect 119270 141148 119308 141204
rect 119364 141148 119374 141204
rect 145366 141148 145404 141204
rect 145460 141148 145470 141204
rect 173012 141148 185052 141204
rect 185108 141148 186396 141204
rect 186452 141148 186462 141204
rect 214582 141148 214620 141204
rect 214676 141148 214686 141204
rect 219286 141148 219324 141204
rect 219380 141148 219390 141204
rect 244598 141148 244636 141204
rect 244692 141148 244702 141204
rect 314598 141148 314636 141204
rect 314692 141148 314702 141204
rect 319190 141148 319228 141204
rect 319284 141148 319294 141204
rect 340946 141148 340956 141204
rect 341012 141148 345324 141204
rect 345380 141148 345390 141204
rect 373426 141148 373436 141204
rect 373492 141148 374556 141204
rect 374612 141148 374622 141204
rect 414082 141148 414092 141204
rect 414148 141148 414652 141204
rect 414708 141148 414718 141204
rect 418338 141148 418348 141204
rect 418404 141148 419244 141204
rect 419300 141148 419310 141204
rect 463708 141148 474124 141204
rect 474180 141148 474190 141204
rect 534566 141148 534604 141204
rect 534660 141148 534670 141204
rect 544646 141148 544684 141204
rect 544740 141148 544750 141204
rect 173012 141092 173068 141148
rect 463708 141092 463764 141148
rect 85026 141036 85036 141092
rect 85092 141036 173068 141092
rect 373874 141036 373884 141092
rect 373940 141036 463764 141092
rect 331762 140924 331772 140980
rect 331828 140924 416332 140980
rect 416388 140924 503916 140980
rect 503972 140924 503982 140980
rect 117506 140812 117516 140868
rect 117572 140812 217420 140868
rect 217476 140812 217486 140868
rect 391906 140812 391916 140868
rect 391972 140812 392252 140868
rect 392308 140812 491596 140868
rect 491652 140812 491662 140868
rect 124338 140700 124348 140756
rect 124404 140700 125468 140756
rect 125524 140700 175420 140756
rect 175476 140700 175486 140756
rect 393362 140700 393372 140756
rect 393428 140700 393932 140756
rect 393988 140700 493388 140756
rect 493444 140700 493454 140756
rect 93314 140588 93324 140644
rect 93380 140588 103964 140644
rect 104020 140588 193340 140644
rect 193396 140588 193406 140644
rect 245382 140588 245420 140644
rect 245476 140588 303212 140644
rect 303268 140588 303996 140644
rect 304052 140588 304062 140644
rect 335010 140588 335020 140644
rect 335076 140588 433468 140644
rect 433524 140588 434812 140644
rect 434868 140588 434878 140644
rect 484754 140588 484764 140644
rect 484820 140588 533820 140644
rect 533876 140588 533886 140644
rect 100818 140476 100828 140532
rect 100884 140476 192780 140532
rect 192836 140476 192846 140532
rect 216402 140476 216412 140532
rect 216468 140476 316428 140532
rect 316484 140476 316494 140532
rect 392466 140476 392476 140532
rect 392532 140476 392812 140532
rect 392868 140476 493052 140532
rect 493108 140476 493118 140532
rect 97682 140364 97692 140420
rect 97748 140364 191996 140420
rect 192052 140364 192062 140420
rect 217410 140364 217420 140420
rect 217476 140364 317436 140420
rect 317492 140364 317502 140420
rect 385746 140364 385756 140420
rect 385812 140364 486332 140420
rect 486388 140364 486398 140420
rect 96450 140252 96460 140308
rect 96516 140252 190988 140308
rect 191044 140252 191054 140308
rect 193330 140252 193340 140308
rect 193396 140252 293356 140308
rect 293412 140252 293422 140308
rect 391010 140252 391020 140308
rect 391076 140252 491372 140308
rect 491428 140252 491438 140308
rect 185714 140140 185724 140196
rect 185780 140140 285740 140196
rect 285796 140140 285806 140196
rect 336018 140140 336028 140196
rect 336084 140140 417452 140196
rect 417508 140140 498988 140196
rect 499044 140140 499054 140196
rect 191986 140028 191996 140084
rect 192052 140028 292012 140084
rect 292068 140028 292078 140084
rect 292786 140028 292796 140084
rect 292852 140028 392812 140084
rect 392868 140028 392878 140084
rect 433794 140028 433804 140084
rect 433860 140028 484764 140084
rect 484820 140028 484830 140084
rect 190978 139916 190988 139972
rect 191044 139916 291004 139972
rect 291060 139916 390572 139972
rect 390628 139916 391020 139972
rect 391076 139916 391086 139972
rect 116722 139804 116732 139860
rect 116788 139804 216412 139860
rect 216468 139804 216478 139860
rect 285730 139804 285740 139860
rect 285796 139804 385756 139860
rect 385812 139804 385822 139860
rect 174178 139692 174188 139748
rect 174244 139692 274204 139748
rect 274260 139692 373884 139748
rect 373940 139692 374220 139748
rect 374276 139692 374286 139748
rect 133746 139580 133756 139636
rect 133812 139580 233772 139636
rect 233828 139580 233838 139636
rect 292002 139580 292012 139636
rect 292068 139580 391916 139636
rect 391972 139580 391982 139636
rect 192770 139468 192780 139524
rect 192836 139468 292796 139524
rect 292852 139468 292862 139524
rect 293346 139468 293356 139524
rect 293412 139468 393372 139524
rect 393428 139468 393438 139524
rect 57138 139356 57148 139412
rect 57204 139356 61180 139412
rect 61236 139356 61246 139412
rect 223346 139356 223356 139412
rect 223412 139356 314188 139412
rect 314132 139300 314188 139356
rect 595560 139300 597000 139496
rect 96898 139244 96908 139300
rect 96964 139244 102508 139300
rect 234994 139244 235004 139300
rect 235060 139244 312508 139300
rect 312564 139244 312574 139300
rect 314132 139244 323596 139300
rect 323652 139244 420028 139300
rect 568642 139244 568652 139300
rect 568708 139272 597000 139300
rect 568708 139244 595672 139272
rect 102452 139188 102508 139244
rect 419972 139188 420028 139244
rect 102452 139132 196700 139188
rect 196756 139132 196766 139188
rect 233986 139132 233996 139188
rect 234052 139132 315420 139188
rect 315476 139132 315486 139188
rect 330866 139132 330876 139188
rect 330932 139132 417676 139188
rect 417732 139132 417742 139188
rect 419972 139132 423612 139188
rect 423668 139132 424172 139188
rect 424228 139132 495404 139188
rect 495460 139132 495470 139188
rect 496636 139132 500668 139188
rect 500724 139132 500734 139188
rect 123330 139020 123340 139076
rect 123396 139020 126028 139076
rect 175410 139020 175420 139076
rect 175476 139020 275436 139076
rect 275492 139020 275502 139076
rect 345314 139020 345324 139076
rect 345380 139020 445564 139076
rect 445620 139020 445630 139076
rect 125972 138964 126028 139020
rect 496636 138964 496692 139132
rect 496850 139020 496860 139076
rect 496916 139020 496926 139076
rect 125972 138908 223356 138964
rect 223412 138908 223422 138964
rect 259522 138908 259532 138964
rect 259588 138908 260428 138964
rect 260484 138908 260494 138964
rect 263778 138908 263788 138964
rect 263844 138908 363804 138964
rect 363860 138908 363870 138964
rect 418114 138908 418124 138964
rect 418180 138908 496692 138964
rect 496860 138852 496916 139020
rect 122658 138796 122668 138852
rect 122724 138796 185612 138852
rect 185668 138796 185678 138852
rect 196914 138796 196924 138852
rect 196980 138796 296828 138852
rect 296884 138796 396844 138852
rect 396900 138796 397292 138852
rect 397348 138796 496916 138852
rect 118178 138684 118188 138740
rect 118244 138684 218204 138740
rect 218260 138684 317772 138740
rect 317828 138684 317838 138740
rect 333778 138684 333788 138740
rect 333844 138684 433804 138740
rect 433860 138684 433870 138740
rect 434914 138684 434924 138740
rect 434980 138684 484876 138740
rect 484932 138684 484942 138740
rect 135426 138572 135436 138628
rect 135492 138572 234780 138628
rect 234836 138572 234846 138628
rect 275314 138572 275324 138628
rect 275380 138572 375228 138628
rect 375284 138572 475244 138628
rect 475300 138572 475310 138628
rect 392 135800 4172 135828
rect -960 135772 4172 135800
rect 4228 135772 4238 135828
rect -960 135576 480 135772
rect 590146 126252 590156 126308
rect 590212 126280 595672 126308
rect 590212 126252 597000 126280
rect 595560 126056 597000 126252
rect -960 121464 480 121688
rect 590594 113036 590604 113092
rect 590660 113064 595672 113092
rect 590660 113036 597000 113064
rect 595560 112840 597000 113036
rect -960 107380 480 107576
rect -960 107352 19292 107380
rect 392 107324 19292 107352
rect 19348 107324 19358 107380
rect 590818 99820 590828 99876
rect 590884 99848 595672 99876
rect 590884 99820 597000 99848
rect 595560 99624 597000 99820
rect -960 93268 480 93464
rect -960 93240 12572 93268
rect 392 93212 12572 93240
rect 12628 93212 12638 93268
rect 590594 86604 590604 86660
rect 590660 86632 595672 86660
rect 590660 86604 597000 86632
rect 595560 86408 597000 86604
rect -960 79128 480 79352
rect 590482 73388 590492 73444
rect 590548 73416 595672 73444
rect 590548 73388 597000 73416
rect 595560 73192 597000 73388
rect 392 65240 7532 65268
rect -960 65212 7532 65240
rect 7588 65212 7598 65268
rect -960 65016 480 65212
rect 595560 60004 597000 60200
rect 566962 59948 566972 60004
rect 567028 59976 597000 60004
rect 567028 59948 595672 59976
rect -960 50932 480 51128
rect -960 50904 14252 50932
rect 392 50876 14252 50904
rect 14308 50876 14318 50932
rect 590482 46956 590492 47012
rect 590548 46984 595672 47012
rect 590548 46956 597000 46984
rect 595560 46760 597000 46956
rect 142818 40236 142828 40292
rect 142884 40236 152012 40292
rect 152068 40236 152078 40292
rect 97010 39452 97020 39508
rect 97076 39452 149772 39508
rect 149828 39452 149838 39508
rect 195906 39452 195916 39508
rect 195972 39452 249228 39508
rect 249284 39452 249294 39508
rect 449474 39452 449484 39508
rect 449540 39452 460684 39508
rect 460740 39452 460750 39508
rect 456194 37996 456204 38052
rect 456260 37996 489244 38052
rect 489300 37996 489310 38052
rect 58706 37884 58716 37940
rect 58772 37884 72268 37940
rect 72324 37884 72334 37940
rect 106530 37884 106540 37940
rect 106596 37884 154588 37940
rect 154644 37884 154654 37940
rect 197922 37884 197932 37940
rect 197988 37884 252140 37940
rect 252196 37884 252206 37940
rect 454514 37884 454524 37940
rect 454580 37884 512092 37940
rect 512148 37884 512158 37940
rect 59714 37772 59724 37828
rect 59780 37772 76076 37828
rect 76132 37772 76142 37828
rect 110338 37772 110348 37828
rect 110404 37772 159740 37828
rect 159796 37772 159806 37828
rect 196018 37772 196028 37828
rect 196084 37772 255724 37828
rect 255780 37772 255790 37828
rect 460114 37772 460124 37828
rect 460180 37772 534940 37828
rect 534996 37772 535006 37828
rect -960 36820 480 37016
rect -960 36792 20972 36820
rect 392 36764 20972 36792
rect 21028 36764 21038 36820
rect 119858 36204 119868 36260
rect 119924 36204 155372 36260
rect 155428 36204 155438 36260
rect 209346 36204 209356 36260
rect 209412 36204 259532 36260
rect 259588 36204 259598 36260
rect 95106 36092 95116 36148
rect 95172 36092 149660 36148
rect 149716 36092 149726 36148
rect 201730 36092 201740 36148
rect 201796 36092 255612 36148
rect 255668 36092 255678 36148
rect 355282 36092 355292 36148
rect 355348 36092 437836 36148
rect 437892 36092 437902 36148
rect 460226 36092 460236 36148
rect 460292 36092 540652 36148
rect 540708 36092 540718 36148
rect 457874 34412 457884 34468
rect 457940 34412 517804 34468
rect 517860 34412 517870 34468
rect 595560 33684 597000 33768
rect 55346 33628 55356 33684
rect 55412 33628 597000 33684
rect 595560 33544 597000 33628
rect 207442 32732 207452 32788
rect 207508 32732 257964 32788
rect 258020 32732 258030 32788
rect 451154 32732 451164 32788
rect 451220 32732 529228 32788
rect 529284 32732 529294 32788
rect 203634 31052 203644 31108
rect 203700 31052 257852 31108
rect 257908 31052 257918 31108
rect 199938 29372 199948 29428
rect 200004 29372 258748 29428
rect 258804 29372 258814 29428
rect 83682 26012 83692 26068
rect 83748 26012 121772 26068
rect 121828 26012 121838 26068
rect 18946 24332 18956 24388
rect 19012 24332 26012 24388
rect 26068 24332 26078 24388
rect 87490 24332 87500 24388
rect 87556 24332 147980 24388
rect 148036 24332 148046 24388
rect 451042 24332 451052 24388
rect 451108 24332 506380 24388
rect 506436 24332 506446 24388
rect -960 22708 480 22904
rect -960 22680 22652 22708
rect 392 22652 22652 22680
rect 22708 22652 22718 22708
rect 595560 20356 597000 20552
rect 353602 20300 353612 20356
rect 353668 20328 597000 20356
rect 353668 20300 595672 20328
rect 284722 17612 284732 17668
rect 284788 17612 426412 17668
rect 426468 17612 426478 17668
rect 91298 15932 91308 15988
rect 91364 15932 138572 15988
rect 138628 15932 138638 15988
rect 291442 15932 291452 15988
rect 291508 15932 420700 15988
rect 420756 15932 420766 15988
rect 176978 14252 176988 14308
rect 177044 14252 227612 14308
rect 227668 14252 227678 14308
rect 260754 14252 260764 14308
rect 260820 14252 273868 14308
rect 273924 14252 273934 14308
rect 298162 14252 298172 14308
rect 298228 14252 392140 14308
rect 392196 14252 392206 14308
rect 20850 13356 20860 13412
rect 20916 13356 27692 13412
rect 27748 13356 27758 13412
rect 104626 12572 104636 12628
rect 104692 12572 153020 12628
rect 153076 12572 153086 12628
rect 184594 12572 184604 12628
rect 184660 12572 237692 12628
rect 237748 12572 237758 12628
rect -960 8596 480 8792
rect -960 8568 15932 8596
rect 392 8540 15932 8568
rect 15988 8540 15998 8596
rect 99026 7644 99036 7700
rect 99092 7644 149548 7700
rect 149604 7644 149614 7700
rect 186722 7644 186732 7700
rect 186788 7644 239372 7700
rect 239428 7644 239438 7700
rect 93426 7532 93436 7588
rect 93492 7532 147868 7588
rect 147924 7532 147934 7588
rect 190530 7532 190540 7588
rect 190596 7532 252028 7588
rect 252084 7532 252094 7588
rect 296482 7532 296492 7588
rect 296548 7532 317884 7588
rect 317940 7532 317950 7588
rect 595560 7140 597000 7336
rect 565282 7084 565292 7140
rect 565348 7112 597000 7140
rect 565348 7084 595672 7112
rect 182914 6076 182924 6132
rect 182980 6076 230972 6132
rect 231028 6076 231038 6132
rect 89618 5964 89628 6020
rect 89684 5964 136892 6020
rect 136948 5964 136958 6020
rect 220994 5964 221004 6020
rect 221060 5964 270508 6020
rect 270564 5964 270574 6020
rect 289762 5964 289772 6020
rect 289828 5964 295036 6020
rect 295092 5964 295102 6020
rect 299842 5964 299852 6020
rect 299908 5964 312172 6020
rect 312228 5964 312238 6020
rect 452834 5964 452844 6020
rect 452900 5964 466396 6020
rect 466452 5964 466462 6020
rect 101042 5852 101052 5908
rect 101108 5852 152908 5908
rect 152964 5852 152974 5908
rect 215282 5852 215292 5908
rect 215348 5852 269388 5908
rect 269444 5852 269454 5908
rect 293122 5852 293132 5908
rect 293188 5852 409276 5908
rect 409332 5852 409342 5908
rect 454402 5852 454412 5908
rect 454468 5852 500668 5908
rect 500724 5852 500734 5908
rect 139122 5068 139132 5124
rect 139188 5068 140252 5124
rect 140308 5068 140318 5124
rect 279682 5068 279692 5124
rect 279748 5068 283612 5124
rect 283668 5068 283678 5124
rect 288082 5068 288092 5124
rect 288148 5068 289324 5124
rect 289380 5068 289390 5124
rect 294802 5068 294812 5124
rect 294868 5068 300748 5124
rect 300804 5068 300814 5124
rect 55346 4956 55356 5012
rect 55412 4956 56252 5012
rect 56308 4956 56318 5012
rect 146738 4956 146748 5012
rect 146804 4956 152124 5012
rect 152180 4956 152190 5012
rect 350466 4956 350476 5012
rect 350532 4956 363580 5012
rect 363636 4956 363646 5012
rect 30594 4844 30604 4900
rect 30660 4844 32732 4900
rect 32788 4844 32798 4900
rect 40114 4844 40124 4900
rect 40180 4844 44492 4900
rect 44548 4844 44558 4900
rect 141026 4844 141036 4900
rect 141092 4844 157276 4900
rect 157332 4844 157342 4900
rect 355282 4844 355292 4900
rect 355348 4844 375004 4900
rect 375060 4844 375070 4900
rect 133410 4732 133420 4788
rect 133476 4732 143612 4788
rect 143668 4732 143678 4788
rect 144834 4732 144844 4788
rect 144900 4732 152012 4788
rect 152068 4732 152078 4788
rect 350242 4732 350252 4788
rect 350308 4732 380716 4788
rect 380772 4732 380782 4788
rect 121986 4620 121996 4676
rect 122052 4620 130172 4676
rect 130228 4620 130238 4676
rect 135314 4620 135324 4676
rect 135380 4620 155372 4676
rect 155428 4620 155438 4676
rect 160850 4620 160860 4676
rect 160916 4620 175084 4676
rect 175140 4620 175150 4676
rect 238130 4620 238140 4676
rect 238196 4620 247772 4676
rect 247828 4620 247838 4676
rect 353602 4620 353612 4676
rect 353668 4620 386428 4676
rect 386484 4620 386494 4676
rect 456082 4620 456092 4676
rect 456148 4620 472108 4676
rect 472164 4620 472174 4676
rect 34514 4508 34524 4564
rect 34580 4508 51212 4564
rect 51268 4508 51278 4564
rect 127586 4508 127596 4564
rect 127652 4508 148876 4564
rect 148932 4508 148942 4564
rect 150668 4508 157500 4564
rect 157556 4508 157566 4564
rect 163874 4508 163884 4564
rect 163940 4508 192332 4564
rect 192388 4508 192398 4564
rect 211474 4508 211484 4564
rect 211540 4508 257852 4564
rect 257908 4508 257918 4564
rect 337652 4508 347900 4564
rect 347956 4508 347966 4564
rect 360322 4508 360332 4564
rect 360388 4508 403564 4564
rect 403620 4508 403630 4564
rect 457762 4508 457772 4564
rect 457828 4508 477820 4564
rect 477876 4508 477886 4564
rect 15362 4396 15372 4452
rect 15428 4396 20188 4452
rect 60162 4396 60172 4452
rect 60228 4396 66556 4452
rect 66612 4396 66622 4452
rect 125794 4396 125804 4452
rect 125860 4396 150444 4452
rect 150500 4396 150510 4452
rect 20132 4340 20188 4396
rect 13346 4284 13356 4340
rect 13412 4284 17612 4340
rect 17668 4284 17678 4340
rect 20132 4284 29372 4340
rect 29428 4284 29438 4340
rect 32498 4284 32508 4340
rect 32564 4284 34412 4340
rect 34468 4284 34478 4340
rect 42018 4284 42028 4340
rect 42084 4284 42812 4340
rect 42868 4284 42878 4340
rect 45724 4284 47852 4340
rect 47908 4284 47918 4340
rect 59938 4284 59948 4340
rect 60004 4284 60844 4340
rect 60900 4284 60910 4340
rect 68674 4284 68684 4340
rect 68740 4284 81452 4340
rect 81508 4284 81518 4340
rect 85810 4284 85820 4340
rect 85876 4284 89852 4340
rect 89908 4284 89918 4340
rect 123890 4284 123900 4340
rect 123956 4284 148652 4340
rect 148708 4284 148718 4340
rect 45724 4228 45780 4284
rect 150668 4228 150724 4508
rect 161970 4396 161980 4452
rect 162036 4396 195692 4452
rect 195748 4396 195758 4452
rect 205762 4396 205772 4452
rect 205828 4396 259532 4452
rect 259588 4396 259598 4452
rect 152450 4284 152460 4340
rect 152516 4284 160412 4340
rect 160468 4284 160478 4340
rect 169586 4284 169596 4340
rect 169652 4284 188972 4340
rect 189028 4284 189038 4340
rect 192434 4284 192444 4340
rect 192500 4284 247548 4340
rect 247604 4284 247614 4340
rect 266690 4284 266700 4340
rect 266756 4284 267036 4340
rect 267092 4284 267102 4340
rect 337652 4228 337708 4508
rect 351922 4396 351932 4452
rect 351988 4396 397852 4452
rect 397908 4396 397918 4452
rect 452722 4396 452732 4452
rect 452788 4396 483532 4452
rect 483588 4396 483598 4452
rect 346658 4284 346668 4340
rect 346724 4284 348012 4340
rect 348068 4284 348078 4340
rect 348562 4284 348572 4340
rect 348628 4284 414988 4340
rect 415044 4284 415054 4340
rect 449362 4284 449372 4340
rect 449428 4284 494956 4340
rect 495012 4284 495022 4340
rect 549332 4284 559468 4340
rect 559524 4284 559534 4340
rect 549332 4228 549388 4284
rect 17266 4172 17276 4228
rect 17332 4172 24332 4228
rect 24388 4172 24398 4228
rect 26786 4172 26796 4228
rect 26852 4172 45780 4228
rect 47730 4172 47740 4228
rect 47796 4172 49532 4228
rect 49588 4172 49598 4228
rect 60274 4172 60284 4228
rect 60340 4172 64652 4228
rect 64708 4172 64718 4228
rect 70326 4172 70364 4228
rect 70420 4172 70430 4228
rect 78194 4172 78204 4228
rect 78260 4172 78876 4228
rect 78932 4172 78942 4228
rect 80098 4172 80108 4228
rect 80164 4172 80556 4228
rect 80612 4172 80622 4228
rect 82002 4172 82012 4228
rect 82068 4172 86492 4228
rect 86548 4172 86558 4228
rect 102946 4172 102956 4228
rect 103012 4172 104972 4228
rect 105028 4172 105038 4228
rect 108658 4172 108668 4228
rect 108724 4172 109116 4228
rect 109172 4172 109182 4228
rect 112438 4172 112476 4228
rect 112532 4172 112542 4228
rect 114370 4172 114380 4228
rect 114436 4172 116732 4228
rect 116788 4172 116798 4228
rect 118178 4172 118188 4228
rect 118244 4172 119196 4228
rect 119252 4172 119262 4228
rect 125972 4172 150724 4228
rect 156146 4172 156156 4228
rect 156212 4172 157052 4228
rect 157108 4172 157118 4228
rect 167878 4172 167916 4228
rect 167972 4172 167982 4228
rect 171266 4172 171276 4228
rect 171332 4172 171388 4228
rect 171444 4172 171454 4228
rect 173012 4172 185612 4228
rect 185668 4172 185678 4228
rect 194338 4172 194348 4228
rect 194404 4172 195916 4228
rect 195972 4172 195982 4228
rect 196532 4172 243628 4228
rect 243842 4172 243852 4228
rect 243908 4172 245196 4228
rect 245252 4172 245262 4228
rect 250338 4172 250348 4228
rect 250404 4172 250414 4228
rect 260306 4172 260316 4228
rect 260372 4172 272188 4228
rect 272244 4172 272254 4228
rect 277862 4172 277900 4228
rect 277956 4172 277966 4228
rect 304882 4172 304892 4228
rect 304948 4172 306460 4228
rect 306516 4172 306526 4228
rect 322578 4172 322588 4228
rect 322644 4172 323596 4228
rect 323652 4172 323662 4228
rect 329270 4172 329308 4228
rect 329364 4172 329374 4228
rect 335234 4172 335244 4228
rect 335300 4172 337708 4228
rect 340946 4172 340956 4228
rect 341012 4172 347788 4228
rect 347844 4172 347854 4228
rect 358642 4172 358652 4228
rect 358708 4172 432124 4228
rect 432180 4172 432190 4228
rect 443762 4172 443772 4228
rect 443828 4172 447468 4228
rect 447524 4172 447534 4228
rect 459442 4172 459452 4228
rect 459508 4172 523516 4228
rect 523572 4172 523582 4228
rect 546578 4172 546588 4228
rect 546644 4172 549388 4228
rect 558002 4172 558012 4228
rect 558068 4172 559580 4228
rect 559636 4172 559646 4228
rect 125972 4116 126028 4172
rect 173012 4116 173068 4172
rect 196532 4116 196588 4172
rect 243572 4116 243628 4172
rect 250348 4116 250404 4172
rect 22978 4060 22988 4116
rect 23044 4060 31052 4116
rect 31108 4060 31118 4116
rect 60050 4060 60060 4116
rect 60116 4060 62748 4116
rect 62804 4060 62814 4116
rect 67172 4060 74172 4116
rect 74228 4060 74238 4116
rect 116274 4060 116284 4116
rect 116340 4060 126028 4116
rect 131506 4060 131516 4116
rect 131572 4060 135212 4116
rect 135268 4060 135278 4116
rect 143602 4060 143612 4116
rect 143668 4060 152572 4116
rect 152628 4060 152638 4116
rect 165778 4060 165788 4116
rect 165844 4060 173068 4116
rect 179106 4060 179116 4116
rect 179172 4060 179676 4116
rect 179732 4060 179742 4116
rect 181010 4060 181020 4116
rect 181076 4060 182252 4116
rect 182308 4060 182318 4116
rect 188626 4060 188636 4116
rect 188692 4060 196588 4116
rect 226678 4060 226716 4116
rect 226772 4060 226782 4116
rect 232418 4060 232428 4116
rect 232484 4060 233436 4116
rect 233492 4060 233502 4116
rect 243572 4060 250404 4116
rect 356962 4060 356972 4116
rect 357028 4060 369292 4116
rect 369348 4060 369358 4116
rect 67172 4004 67228 4060
rect 58594 3948 58604 4004
rect 58660 3948 67228 4004
rect 129602 3948 129612 4004
rect 129668 3948 133532 4004
rect 133588 3948 133598 4004
rect 173394 3836 173404 3892
rect 173460 3836 180572 3892
rect 180628 3836 180638 3892
rect 137190 3388 137228 3444
rect 137284 3388 137294 3444
<< via3 >>
rect 584668 591276 584724 591332
rect 51996 588588 52052 588644
rect 50316 575372 50372 575428
rect 4172 558908 4228 558964
rect 212492 554316 212548 554372
rect 301084 550060 301140 550116
rect 301756 549948 301812 550004
rect 301868 549836 301924 549892
rect 387212 549724 387268 549780
rect 362572 549500 362628 549556
rect 323148 549388 323204 549444
rect 328076 549388 328132 549444
rect 333004 549388 333060 549444
rect 337932 549388 337988 549444
rect 342860 549388 342916 549444
rect 347788 549388 347844 549444
rect 352716 549388 352772 549444
rect 357644 549388 357700 549444
rect 392140 549388 392196 549444
rect 386988 549164 387044 549220
rect 392140 549164 392196 549220
rect 431676 549164 431732 549220
rect 333004 549052 333060 549108
rect 303436 548940 303492 548996
rect 342860 548940 342916 548996
rect 468300 548940 468356 548996
rect 590156 548940 590212 548996
rect 300860 548828 300916 548884
rect 352716 548828 352772 548884
rect 468524 548828 468580 548884
rect 386988 548716 387044 548772
rect 387212 548716 387268 548772
rect 431676 548716 431732 548772
rect 446012 548716 446068 548772
rect 301644 548492 301700 548548
rect 362572 548492 362628 548548
rect 303212 548380 303268 548436
rect 337932 548380 337988 548436
rect 357644 548380 357700 548436
rect 467628 548380 467684 548436
rect 323148 548268 323204 548324
rect 300972 547148 301028 547204
rect 323148 547148 323204 547204
rect 301532 547036 301588 547092
rect 357644 547036 357700 547092
rect 300748 546924 300804 546980
rect 328076 546924 328132 546980
rect 303324 546812 303380 546868
rect 347788 546812 347844 546868
rect 468188 546812 468244 546868
rect 4284 545020 4340 545076
rect 548156 537740 548212 537796
rect 549388 535948 549444 536004
rect 590604 535836 590660 535892
rect 529340 534268 529396 534324
rect 529340 533372 529396 533428
rect 549500 533372 549556 533428
rect 4172 530796 4228 530852
rect 556220 529340 556276 529396
rect 590492 522732 590548 522788
rect 300524 521724 300580 521780
rect 300636 520268 300692 520324
rect 556108 518812 556164 518868
rect 300524 516796 300580 516852
rect 300636 513548 300692 513604
rect 300860 511196 300916 511252
rect 590716 509292 590772 509348
rect 300748 505820 300804 505876
rect 300972 503132 301028 503188
rect 176988 501676 177044 501732
rect 171500 501564 171556 501620
rect 176988 500556 177044 500612
rect 171500 499996 171556 500052
rect 301084 497196 301140 497252
rect 590492 496076 590548 496132
rect 467628 495516 467684 495572
rect 468636 489468 468692 489524
rect 468188 483420 468244 483476
rect 468300 477372 468356 477428
rect 63756 476252 63812 476308
rect 467852 471324 467908 471380
rect 590828 469644 590884 469700
rect 590604 456428 590660 456484
rect 554428 455196 554484 455252
rect 293132 452732 293188 452788
rect 533036 451500 533092 451556
rect 481628 451388 481684 451444
rect 481404 451276 481460 451332
rect 481516 451164 481572 451220
rect 481292 451052 481348 451108
rect 478268 450604 478324 450660
rect 590828 450604 590884 450660
rect 474908 450492 474964 450548
rect 478492 450492 478548 450548
rect 480508 450380 480564 450436
rect 554428 450380 554484 450436
rect 468636 450268 468692 450324
rect 480620 450268 480676 450324
rect 533036 450156 533092 450212
rect 526652 448476 526708 448532
rect 521612 447356 521668 447412
rect 288092 437612 288148 437668
rect 298396 436156 298452 436212
rect 164556 433356 164612 433412
rect 166236 433356 166292 433412
rect 169596 433356 169652 433412
rect 267036 433356 267092 433412
rect 268716 433356 268772 433412
rect 300748 432908 300804 432964
rect 212492 432684 212548 432740
rect 121996 432572 122052 432628
rect 457772 432572 457828 432628
rect 512316 432572 512372 432628
rect 474572 432236 474628 432292
rect 482972 432124 483028 432180
rect 498876 432124 498932 432180
rect 76412 432012 76468 432068
rect 276444 432012 276500 432068
rect 502908 432012 502964 432068
rect 4956 431900 5012 431956
rect 82908 431900 82964 431956
rect 519036 431900 519092 431956
rect 77532 431788 77588 431844
rect 483084 431788 483140 431844
rect 523068 431788 523124 431844
rect 300860 431004 300916 431060
rect 301084 430892 301140 430948
rect 288092 430668 288148 430724
rect 278012 430556 278068 430612
rect 298284 430444 298340 430500
rect 293244 430332 293300 430388
rect 69468 430220 69524 430276
rect 298620 430220 298676 430276
rect 464604 430220 464660 430276
rect 294924 430108 294980 430164
rect 590828 430108 590884 430164
rect 66668 429996 66724 430052
rect 212492 429996 212548 430052
rect 278124 429996 278180 430052
rect 56476 429884 56532 429940
rect 300972 429884 301028 429940
rect 478380 429884 478436 429940
rect 298732 429548 298788 429604
rect 291564 429436 291620 429492
rect 478156 429436 478212 429492
rect 74844 429324 74900 429380
rect 461132 429324 461188 429380
rect 249564 429212 249620 429268
rect 252252 429212 252308 429268
rect 260316 429212 260372 429268
rect 263676 429212 263732 429268
rect 289884 429212 289940 429268
rect 464492 429212 464548 429268
rect 279692 429100 279748 429156
rect 60620 428540 60676 428596
rect 83244 428428 83300 428484
rect 298956 428428 299012 428484
rect 252252 427756 252308 427812
rect 301084 427756 301140 427812
rect 249564 427644 249620 427700
rect 83580 427532 83636 427588
rect 295260 427532 295316 427588
rect 83356 427420 83412 427476
rect 295036 427420 295092 427476
rect 284956 427308 285012 427364
rect 296492 427196 296548 427252
rect 56364 427084 56420 427140
rect 300860 427084 300916 427140
rect 590716 416780 590772 416836
rect 56588 413644 56644 413700
rect 57036 412300 57092 412356
rect 451052 411852 451108 411908
rect 449372 410284 449428 410340
rect 60172 409164 60228 409220
rect 456092 408716 456148 408772
rect 60284 407708 60340 407764
rect 452732 407148 452788 407204
rect 474796 405580 474852 405636
rect 60508 404684 60564 404740
rect 454412 404012 454468 404068
rect 4284 403900 4340 403956
rect 591052 403564 591108 403620
rect 468636 403340 468692 403396
rect 480620 403116 480676 403172
rect 301756 402668 301812 402724
rect 472892 402444 472948 402500
rect 300748 402332 300804 402388
rect 478380 401212 478436 401268
rect 480508 401100 480564 401156
rect 474684 400876 474740 400932
rect 301644 400652 301700 400708
rect 480508 400652 480564 400708
rect 301532 400540 301588 400596
rect 480620 400540 480676 400596
rect 298060 399644 298116 399700
rect 298508 399532 298564 399588
rect 478044 399532 478100 399588
rect 549500 399532 549556 399588
rect 298956 399420 299012 399476
rect 478268 399420 478324 399476
rect 298172 397964 298228 398020
rect 478156 397964 478212 398020
rect 549388 394156 549444 394212
rect 56700 392140 56756 392196
rect 56812 390796 56868 390852
rect 273196 390572 273252 390628
rect 474796 390572 474852 390628
rect 548156 390572 548212 390628
rect 590940 390348 590996 390404
rect 56476 389452 56532 389508
rect 273532 388780 273588 388836
rect 56924 388108 56980 388164
rect 451052 387436 451108 387492
rect 56364 386764 56420 386820
rect 449372 386092 449428 386148
rect 56140 385420 56196 385476
rect 456092 384748 456148 384804
rect 273644 383964 273700 384020
rect 472892 383964 472948 384020
rect 452732 383404 452788 383460
rect 60284 383292 60340 383348
rect 53676 382732 53732 382788
rect 273196 382060 273252 382116
rect 484764 381836 484820 381892
rect 54348 381388 54404 381444
rect 454412 380716 454468 380772
rect 484764 380716 484820 380772
rect 273756 380604 273812 380660
rect 474684 380604 474740 380660
rect 300972 380380 301028 380436
rect 525868 380380 525924 380436
rect 57932 380044 57988 380100
rect 459452 379932 459508 379988
rect 273644 379372 273700 379428
rect 276332 378812 276388 378868
rect 53564 378700 53620 378756
rect 273756 378028 273812 378084
rect 494844 377916 494900 377972
rect 498876 377916 498932 377972
rect 521052 377916 521108 377972
rect 521612 377916 521668 377972
rect 478156 377468 478212 377524
rect 56812 377356 56868 377412
rect 590156 377132 590212 377188
rect 60172 375340 60228 375396
rect 60732 374668 60788 374724
rect 56700 373324 56756 373380
rect 56588 371980 56644 372036
rect 273756 371308 273812 371364
rect 60172 368620 60228 368676
rect 273756 368620 273812 368676
rect 60732 367948 60788 368004
rect 273756 367276 273812 367332
rect 60732 366604 60788 366660
rect 273756 365932 273812 365988
rect 58492 365260 58548 365316
rect 273756 364588 273812 364644
rect 60060 363916 60116 363972
rect 273084 363244 273140 363300
rect 56476 362572 56532 362628
rect 273756 361900 273812 361956
rect 4172 361564 4228 361620
rect 55020 361228 55076 361284
rect 273756 360556 273812 360612
rect 56364 359884 56420 359940
rect 273308 359212 273364 359268
rect 54796 358540 54852 358596
rect 273644 357868 273700 357924
rect 53452 357196 53508 357252
rect 273756 356524 273812 356580
rect 53228 355852 53284 355908
rect 273756 355180 273812 355236
rect 53340 354508 53396 354564
rect 56252 353164 56308 353220
rect 54908 351820 54964 351876
rect 273644 351148 273700 351204
rect 591052 350700 591108 350756
rect 60508 350028 60564 350084
rect 273756 349804 273812 349860
rect 54684 349132 54740 349188
rect 521612 348572 521668 348628
rect 273756 348460 273812 348516
rect 54572 347788 54628 347844
rect 4172 347452 4228 347508
rect 284732 347116 284788 347172
rect 60284 346444 60340 346500
rect 291452 345772 291508 345828
rect 498988 345324 499044 345380
rect 502348 345324 502404 345380
rect 505708 345324 505764 345380
rect 495964 344876 496020 344932
rect 479948 344652 480004 344708
rect 479724 344540 479780 344596
rect 60508 344428 60564 344484
rect 272972 344428 273028 344484
rect 480172 344428 480228 344484
rect 509404 344428 509460 344484
rect 512764 344428 512820 344484
rect 516124 344428 516180 344484
rect 519484 344428 519540 344484
rect 293132 343084 293188 343140
rect 273196 341740 273252 341796
rect 273756 340396 273812 340452
rect 298172 339052 298228 339108
rect 51996 338380 52052 338436
rect 475468 338380 475524 338436
rect 273308 337708 273364 337764
rect 475468 337484 475524 337540
rect 591164 337484 591220 337540
rect 58716 337036 58772 337092
rect 475580 336588 475636 336644
rect 273084 336364 273140 336420
rect 60732 335692 60788 335748
rect 475468 335692 475524 335748
rect 60172 335020 60228 335076
rect 4172 333116 4228 333172
rect 60508 333004 60564 333060
rect 475468 333004 475524 333060
rect 475468 332108 475524 332164
rect 53116 331660 53172 331716
rect 475580 331212 475636 331268
rect 475468 330316 475524 330372
rect 60172 329420 60228 329476
rect 475692 329420 475748 329476
rect 58156 328972 58212 329028
rect 390572 328524 390628 328580
rect 60732 327628 60788 327684
rect 476252 327628 476308 327684
rect 475468 326732 475524 326788
rect 58268 326284 58324 326340
rect 60396 324268 60452 324324
rect 58044 323596 58100 323652
rect 55244 322252 55300 322308
rect 296492 321580 296548 321636
rect 475468 321356 475524 321412
rect 58380 320908 58436 320964
rect 472892 320460 472948 320516
rect 299852 320236 299908 320292
rect 54460 319564 54516 319620
rect 473116 319564 473172 319620
rect 4284 319004 4340 319060
rect 475580 318668 475636 318724
rect 475468 317772 475524 317828
rect 294812 317548 294868 317604
rect 289772 316204 289828 316260
rect 475468 315084 475524 315140
rect 288092 314860 288148 314916
rect 279692 313516 279748 313572
rect 475468 313292 475524 313348
rect 50316 312844 50372 312900
rect 277676 312172 277732 312228
rect 55356 311500 55412 311556
rect 476588 311500 476644 311556
rect 591276 311052 591332 311108
rect 272188 310828 272244 310884
rect 476924 310604 476980 310660
rect 58716 310156 58772 310212
rect 476364 309708 476420 309764
rect 58604 308812 58660 308868
rect 475468 308812 475524 308868
rect 273868 308140 273924 308196
rect 476252 307916 476308 307972
rect 60732 307468 60788 307524
rect 476700 307020 476756 307076
rect 57036 306124 57092 306180
rect 476476 306124 476532 306180
rect 476140 305228 476196 305284
rect 4396 304892 4452 304948
rect 60284 304780 60340 304836
rect 476812 304332 476868 304388
rect 55132 303436 55188 303492
rect 477036 303436 477092 303492
rect 388108 302316 388164 302372
rect 56028 302092 56084 302148
rect 55356 300860 55412 300916
rect 54460 300748 54516 300804
rect 57036 300748 57092 300804
rect 388108 300636 388164 300692
rect 388220 300524 388276 300580
rect 270508 298732 270564 298788
rect 590828 297836 590884 297892
rect 269388 297388 269444 297444
rect 388220 297276 388276 297332
rect 388444 297164 388500 297220
rect 60508 296716 60564 296772
rect 56924 295372 56980 295428
rect 476140 293916 476196 293972
rect 56140 292684 56196 292740
rect 288316 292684 288372 292740
rect 56476 292236 56532 292292
rect 293244 292236 293300 292292
rect 388108 292236 388164 292292
rect 56588 292124 56644 292180
rect 289884 292124 289940 292180
rect 56812 292012 56868 292068
rect 283052 292012 283108 292068
rect 56364 291900 56420 291956
rect 281372 291900 281428 291956
rect 278236 291788 278292 291844
rect 56252 291676 56308 291732
rect 276332 291676 276388 291732
rect 56700 291564 56756 291620
rect 274652 291564 274708 291620
rect 247772 291452 247828 291508
rect 4956 290780 5012 290836
rect 388108 290556 388164 290612
rect 63756 290108 63812 290164
rect 245196 289772 245252 289828
rect 475468 288988 475524 289044
rect 180572 286972 180628 287028
rect 155372 286860 155428 286916
rect 177212 286860 177268 286916
rect 167132 286748 167188 286804
rect 152012 286636 152068 286692
rect 121772 286524 121828 286580
rect 149660 286524 149716 286580
rect 168812 286524 168868 286580
rect 140252 286412 140308 286468
rect 200732 286412 200788 286468
rect 230972 286412 231028 286468
rect 258748 286412 258804 286468
rect 123452 286300 123508 286356
rect 147980 286300 148036 286356
rect 255724 286300 255780 286356
rect 136892 286188 136948 286244
rect 149548 286188 149604 286244
rect 149772 285964 149828 286020
rect 257964 285852 258020 285908
rect 152908 285740 152964 285796
rect 197372 285740 197428 285796
rect 227612 285740 227668 285796
rect 252028 285740 252084 285796
rect 259532 285740 259588 285796
rect 124348 285628 124404 285684
rect 138572 285628 138628 285684
rect 147868 285628 147924 285684
rect 153020 285628 153076 285684
rect 154588 285628 154644 285684
rect 159740 285628 159796 285684
rect 164668 285628 164724 285684
rect 173068 285628 173124 285684
rect 174748 285628 174804 285684
rect 178108 285628 178164 285684
rect 183148 285628 183204 285684
rect 184828 285628 184884 285684
rect 188188 285628 188244 285684
rect 191548 285628 191604 285684
rect 194908 285628 194964 285684
rect 198268 285628 198324 285684
rect 203308 285628 203364 285684
rect 208348 285628 208404 285684
rect 213388 285628 213444 285684
rect 215068 285628 215124 285684
rect 218428 285628 218484 285684
rect 221788 285628 221844 285684
rect 225148 285628 225204 285684
rect 228508 285628 228564 285684
rect 231868 285628 231924 285684
rect 237692 285628 237748 285684
rect 239372 285628 239428 285684
rect 243516 285628 243572 285684
rect 246876 285628 246932 285684
rect 249228 285628 249284 285684
rect 252140 285628 252196 285684
rect 255612 285628 255668 285684
rect 257852 285628 257908 285684
rect 260428 285628 260484 285684
rect 265468 285628 265524 285684
rect 104972 285068 105028 285124
rect 590156 284844 590212 284900
rect 116732 283276 116788 283332
rect 81452 281372 81508 281428
rect 171276 281372 171332 281428
rect 54908 281036 54964 281092
rect 476252 281036 476308 281092
rect 54684 280700 54740 280756
rect 476476 280700 476532 280756
rect 83132 280476 83188 280532
rect 473116 280476 473172 280532
rect 83356 280364 83412 280420
rect 472892 280364 472948 280420
rect 304892 279916 304948 279972
rect 60620 278236 60676 278292
rect 58268 278012 58324 278068
rect 590828 278012 590884 278068
rect 58380 272972 58436 273028
rect 590492 272972 590548 273028
rect 74732 271404 74788 271460
rect 56924 271292 56980 271348
rect 566972 271292 567028 271348
rect 479612 269724 479668 269780
rect 288204 268044 288260 268100
rect 56028 267932 56084 267988
rect 572012 267932 572068 267988
rect 477932 264684 477988 264740
rect 76412 264572 76468 264628
rect 55356 261212 55412 261268
rect 590716 261212 590772 261268
rect 73052 259532 73108 259588
rect 590604 259532 590660 259588
rect 364252 259084 364308 259140
rect 375004 259084 375060 259140
rect 385756 259084 385812 259140
rect 390572 259084 390628 259140
rect 393932 259084 393988 259140
rect 397292 259084 397348 259140
rect 373884 258972 373940 259028
rect 392252 258972 392308 259028
rect 392476 258972 392532 259028
rect 385420 258860 385476 258916
rect 412412 258748 412468 258804
rect 414092 258748 414148 258804
rect 424396 258748 424452 258804
rect 363916 258636 363972 258692
rect 373772 258636 373828 258692
rect 374892 258636 374948 258692
rect 433468 258636 433524 258692
rect 434252 258524 434308 258580
rect 424060 258412 424116 258468
rect 434140 258412 434196 258468
rect 434588 258412 434644 258468
rect 444668 258412 444724 258468
rect 445340 258412 445396 258468
rect 572012 258188 572068 258244
rect 86492 257964 86548 258020
rect 4172 248444 4228 248500
rect 4172 234556 4228 234612
rect 590828 231980 590884 232036
rect 89852 231084 89908 231140
rect 133532 230972 133588 231028
rect 70364 227724 70420 227780
rect 109116 222572 109172 222628
rect 590716 218764 590772 218820
rect 66668 213276 66724 213332
rect 130172 212716 130228 212772
rect 135212 210924 135268 210980
rect 119196 210812 119252 210868
rect 182252 210812 182308 210868
rect 62972 209916 63028 209972
rect 112476 209356 112532 209412
rect 4172 206332 4228 206388
rect 590156 205548 590212 205604
rect 590604 192332 590660 192388
rect 329308 163772 329364 163828
rect 322588 162092 322644 162148
rect 60508 160524 60564 160580
rect 590828 160524 590884 160580
rect 233436 160300 233492 160356
rect 267036 160188 267092 160244
rect 226716 158956 226772 159012
rect 80556 158844 80612 158900
rect 123452 158844 123508 158900
rect 191548 158844 191604 158900
rect 78876 158732 78932 158788
rect 124348 158732 124404 158788
rect 179676 158732 179732 158788
rect 231868 158732 231924 158788
rect 184828 157052 184884 157108
rect 474572 156268 474628 156324
rect 144508 155484 144564 155540
rect 58044 152460 58100 152516
rect 228508 152348 228564 152404
rect 144732 152124 144788 152180
rect 265468 151116 265524 151172
rect 155484 150556 155540 150612
rect 188188 150556 188244 150612
rect 272188 148764 272244 148820
rect 180572 148652 180628 148708
rect 197372 147196 197428 147252
rect 164668 147084 164724 147140
rect 246876 146188 246932 146244
rect 174748 145740 174804 145796
rect 168812 145628 168868 145684
rect 114716 145516 114772 145572
rect 194908 145404 194964 145460
rect 55244 145292 55300 145348
rect 590604 145292 590660 145348
rect 167132 144172 167188 144228
rect 173068 143948 173124 144004
rect 178108 143836 178164 143892
rect 243516 143836 243572 143892
rect 183148 143724 183204 143780
rect 177212 143612 177268 143668
rect 180572 143612 180628 143668
rect 225148 143612 225204 143668
rect 498988 142828 499044 142884
rect 144732 142716 144788 142772
rect 304780 142716 304836 142772
rect 330876 142716 330932 142772
rect 333452 142716 333508 142772
rect 412412 142716 412468 142772
rect 385532 142604 385588 142660
rect 375116 142492 375172 142548
rect 144508 142380 144564 142436
rect 433692 142380 433748 142436
rect 84924 142268 84980 142324
rect 130956 142268 131012 142324
rect 364252 142268 364308 142324
rect 344652 142044 344708 142100
rect 62188 141932 62244 141988
rect 433692 141932 433748 141988
rect 444668 141932 444724 141988
rect 471996 141932 472052 141988
rect 363692 141820 363748 141876
rect 375116 141820 375172 141876
rect 424396 141820 424452 141876
rect 434364 141708 434420 141764
rect 434588 141708 434644 141764
rect 484428 141708 484484 141764
rect 373436 141596 373492 141652
rect 434588 141484 434644 141540
rect 505596 141484 505652 141540
rect 374780 141372 374836 141428
rect 164444 141260 164500 141316
rect 385532 141260 385588 141316
rect 63756 141148 63812 141204
rect 114716 141148 114772 141204
rect 119308 141148 119364 141204
rect 145404 141148 145460 141204
rect 214620 141148 214676 141204
rect 219324 141148 219380 141204
rect 244636 141148 244692 141204
rect 314636 141148 314692 141204
rect 319228 141148 319284 141204
rect 340956 141148 341012 141204
rect 373436 141148 373492 141204
rect 414092 141148 414148 141204
rect 414652 141148 414708 141204
rect 418348 141148 418404 141204
rect 534604 141148 534660 141204
rect 544684 141148 544740 141204
rect 373884 141036 373940 141092
rect 392252 140812 392308 140868
rect 393932 140700 393988 140756
rect 245420 140588 245476 140644
rect 303996 140588 304052 140644
rect 433468 140588 433524 140644
rect 392476 140476 392532 140532
rect 385756 140364 385812 140420
rect 390572 139916 390628 139972
rect 385756 139804 385812 139860
rect 373884 139692 373940 139748
rect 424172 139132 424228 139188
rect 445564 139020 445620 139076
rect 260428 138908 260484 138964
rect 397292 138796 397348 138852
rect 590156 126252 590212 126308
rect 590604 113036 590660 113092
rect 590828 99820 590884 99876
rect 590492 73388 590548 73444
rect 566972 59948 567028 60004
rect 152012 40236 152068 40292
rect 149772 39452 149828 39508
rect 249228 39452 249284 39508
rect 449484 39452 449540 39508
rect 456204 37996 456260 38052
rect 154588 37884 154644 37940
rect 252140 37884 252196 37940
rect 454524 37884 454580 37940
rect 159740 37772 159796 37828
rect 255724 37772 255780 37828
rect 155372 36204 155428 36260
rect 259532 36204 259588 36260
rect 149660 36092 149716 36148
rect 255612 36092 255668 36148
rect 355292 36092 355348 36148
rect 457884 34412 457940 34468
rect 257964 32732 258020 32788
rect 451164 32732 451220 32788
rect 257852 31052 257908 31108
rect 258748 29372 258804 29428
rect 121772 26012 121828 26068
rect 147980 24332 148036 24388
rect 451052 24332 451108 24388
rect 284732 17612 284788 17668
rect 138572 15932 138628 15988
rect 291452 15932 291508 15988
rect 227612 14252 227668 14308
rect 273868 14252 273924 14308
rect 298172 14252 298228 14308
rect 153020 12572 153076 12628
rect 237692 12572 237748 12628
rect 149548 7644 149604 7700
rect 239372 7644 239428 7700
rect 147868 7532 147924 7588
rect 252028 7532 252084 7588
rect 296492 7532 296548 7588
rect 230972 6076 231028 6132
rect 136892 5964 136948 6020
rect 270508 5964 270564 6020
rect 289772 5964 289828 6020
rect 299852 5964 299908 6020
rect 452844 5964 452900 6020
rect 152908 5852 152964 5908
rect 269388 5852 269444 5908
rect 293132 5852 293188 5908
rect 454412 5852 454468 5908
rect 140252 5068 140308 5124
rect 279692 5068 279748 5124
rect 288092 5068 288148 5124
rect 294812 5068 294868 5124
rect 152124 4956 152180 5012
rect 143612 4732 143668 4788
rect 350252 4732 350308 4788
rect 130172 4620 130228 4676
rect 247772 4620 247828 4676
rect 353612 4620 353668 4676
rect 456092 4620 456148 4676
rect 192332 4508 192388 4564
rect 360332 4508 360388 4564
rect 457772 4508 457828 4564
rect 81452 4284 81508 4340
rect 89852 4284 89908 4340
rect 195692 4396 195748 4452
rect 160412 4284 160468 4340
rect 188972 4284 189028 4340
rect 267036 4284 267092 4340
rect 351932 4396 351988 4452
rect 452732 4396 452788 4452
rect 348572 4284 348628 4340
rect 449372 4284 449428 4340
rect 70364 4172 70420 4228
rect 78876 4172 78932 4228
rect 80556 4172 80612 4228
rect 86492 4172 86548 4228
rect 104972 4172 105028 4228
rect 109116 4172 109172 4228
rect 112476 4172 112532 4228
rect 116732 4172 116788 4228
rect 119196 4172 119252 4228
rect 157052 4172 157108 4228
rect 167916 4172 167972 4228
rect 171276 4172 171332 4228
rect 185612 4172 185668 4228
rect 245196 4172 245252 4228
rect 277900 4172 277956 4228
rect 304892 4172 304948 4228
rect 322588 4172 322644 4228
rect 329308 4172 329364 4228
rect 358652 4172 358708 4228
rect 447468 4172 447524 4228
rect 135212 4060 135268 4116
rect 143612 4060 143668 4116
rect 179676 4060 179732 4116
rect 182252 4060 182308 4116
rect 226716 4060 226772 4116
rect 233436 4060 233492 4116
rect 133532 3948 133588 4004
rect 180572 3836 180628 3892
rect 137228 3388 137284 3444
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 5418 562350 6038 579922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect 4172 558964 4228 558974
rect 4172 557938 4228 558908
rect 4172 557872 4228 557882
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect 4172 551278 4228 551288
rect 4172 530852 4228 551222
rect 4284 548218 4340 548228
rect 4284 545076 4340 548162
rect 4284 545010 4340 545020
rect 4172 530786 4228 530796
rect 5418 544350 6038 561922
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 5418 472350 6038 489922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect 5418 454350 6038 471922
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 4956 431956 5012 431966
rect 4956 430858 5012 431900
rect 4956 430792 5012 430802
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect 4172 430138 4228 430148
rect 4172 361620 4228 430082
rect 4284 426898 4340 426908
rect 4284 403956 4340 426842
rect 4284 403890 4340 403900
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect 4172 361554 4228 361564
rect 5418 400350 6038 417922
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect 5418 382350 6038 399922
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 5418 364350 6038 381922
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect 4172 347698 4228 347708
rect 4172 347508 4228 347642
rect 4172 347442 4228 347452
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect 5418 346350 6038 363922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect 4172 333172 4228 333182
rect 4172 300538 4228 333116
rect 5418 328350 6038 345922
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect 4172 300472 4228 300482
rect 4284 319060 4340 319070
rect 4284 293878 4340 319004
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect 4284 293812 4340 293822
rect 4396 304948 4452 304958
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect 4396 288658 4452 304892
rect 5418 292350 6038 309922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 4396 288592 4452 288602
rect 4956 290836 5012 290846
rect 4956 283798 5012 290780
rect 4956 283732 5012 283742
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect 5418 274350 6038 291922
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect 5418 256350 6038 273922
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 4172 248518 4228 248538
rect 4172 248434 4228 248444
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 4172 235198 4228 235208
rect 4172 234612 4228 235142
rect 4172 234546 4228 234556
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 4172 206578 4228 206588
rect 4172 206388 4228 206522
rect 4172 206322 4228 206332
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 5418 148350 6038 165922
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect 5418 4350 6038 21922
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 568350 9758 585922
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 9138 532350 9758 549922
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 9138 478350 9758 495922
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 9138 406350 9758 423922
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 9138 370350 9758 387922
rect 9138 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 9758 370350
rect 9138 370226 9758 370294
rect 9138 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 9758 370226
rect 9138 370102 9758 370170
rect 9138 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 9758 370102
rect 9138 369978 9758 370046
rect 9138 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 9758 369978
rect 9138 352350 9758 369922
rect 9138 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 9758 352350
rect 9138 352226 9758 352294
rect 9138 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 9758 352226
rect 9138 352102 9758 352170
rect 9138 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 9758 352102
rect 9138 351978 9758 352046
rect 9138 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 9758 351978
rect 9138 334350 9758 351922
rect 9138 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 9758 334350
rect 9138 334226 9758 334294
rect 9138 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 9758 334226
rect 9138 334102 9758 334170
rect 9138 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 9758 334102
rect 9138 333978 9758 334046
rect 9138 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 9758 333978
rect 9138 316350 9758 333922
rect 9138 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 9758 316350
rect 9138 316226 9758 316294
rect 9138 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 9758 316226
rect 9138 316102 9758 316170
rect 9138 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 9758 316102
rect 9138 315978 9758 316046
rect 9138 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 9758 315978
rect 9138 298350 9758 315922
rect 9138 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 9758 298350
rect 9138 298226 9758 298294
rect 9138 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 9758 298226
rect 9138 298102 9758 298170
rect 9138 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 9758 298102
rect 9138 297978 9758 298046
rect 9138 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 9758 297978
rect 9138 280350 9758 297922
rect 9138 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 9758 280350
rect 9138 280226 9758 280294
rect 9138 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 9758 280226
rect 9138 280102 9758 280170
rect 9138 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 9758 280102
rect 9138 279978 9758 280046
rect 9138 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 9758 279978
rect 9138 262350 9758 279922
rect 9138 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 9758 262350
rect 9138 262226 9758 262294
rect 9138 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 9758 262226
rect 9138 262102 9758 262170
rect 9138 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 9758 262102
rect 9138 261978 9758 262046
rect 9138 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 9758 261978
rect 9138 244350 9758 261922
rect 9138 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 9758 244350
rect 9138 244226 9758 244294
rect 9138 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 9758 244226
rect 9138 244102 9758 244170
rect 9138 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 9758 244102
rect 9138 243978 9758 244046
rect 9138 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 9758 243978
rect 9138 226350 9758 243922
rect 9138 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 9758 226350
rect 9138 226226 9758 226294
rect 9138 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 9758 226226
rect 9138 226102 9758 226170
rect 9138 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 9758 226102
rect 9138 225978 9758 226046
rect 9138 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 9758 225978
rect 9138 208350 9758 225922
rect 9138 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 9758 208350
rect 9138 208226 9758 208294
rect 9138 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 9758 208226
rect 9138 208102 9758 208170
rect 9138 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 9758 208102
rect 9138 207978 9758 208046
rect 9138 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 9758 207978
rect 9138 190350 9758 207922
rect 9138 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 9758 190350
rect 9138 190226 9758 190294
rect 9138 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 9758 190226
rect 9138 190102 9758 190170
rect 9138 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 9758 190102
rect 9138 189978 9758 190046
rect 9138 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 9758 189978
rect 9138 172350 9758 189922
rect 9138 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 9758 172350
rect 9138 172226 9758 172294
rect 9138 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 9758 172226
rect 9138 172102 9758 172170
rect 9138 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 9758 172102
rect 9138 171978 9758 172046
rect 9138 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 9758 171978
rect 9138 154350 9758 171922
rect 9138 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 9758 154350
rect 9138 154226 9758 154294
rect 9138 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 9758 154226
rect 9138 154102 9758 154170
rect 9138 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 9758 154102
rect 9138 153978 9758 154046
rect 9138 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 9758 153978
rect 9138 136350 9758 153922
rect 9138 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 9758 136350
rect 9138 136226 9758 136294
rect 9138 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 9758 136226
rect 9138 136102 9758 136170
rect 9138 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 9758 136102
rect 9138 135978 9758 136046
rect 9138 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 9758 135978
rect 9138 118350 9758 135922
rect 9138 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 9758 118350
rect 9138 118226 9758 118294
rect 9138 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 9758 118226
rect 9138 118102 9758 118170
rect 9138 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 9758 118102
rect 9138 117978 9758 118046
rect 9138 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 9758 117978
rect 9138 100350 9758 117922
rect 9138 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 9758 100350
rect 9138 100226 9758 100294
rect 9138 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 9758 100226
rect 9138 100102 9758 100170
rect 9138 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 9758 100102
rect 9138 99978 9758 100046
rect 9138 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 9758 99978
rect 9138 82350 9758 99922
rect 9138 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 9758 82350
rect 9138 82226 9758 82294
rect 9138 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 9758 82226
rect 9138 82102 9758 82170
rect 9138 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 9758 82102
rect 9138 81978 9758 82046
rect 9138 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 9758 81978
rect 9138 64350 9758 81922
rect 9138 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 9758 64350
rect 9138 64226 9758 64294
rect 9138 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 9758 64226
rect 9138 64102 9758 64170
rect 9138 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 9758 64102
rect 9138 63978 9758 64046
rect 9138 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 9758 63978
rect 9138 46350 9758 63922
rect 9138 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 9758 46350
rect 9138 46226 9758 46294
rect 9138 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 9758 46226
rect 9138 46102 9758 46170
rect 9138 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 9758 46102
rect 9138 45978 9758 46046
rect 9138 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 9758 45978
rect 9138 28350 9758 45922
rect 9138 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 9758 28350
rect 9138 28226 9758 28294
rect 9138 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 9758 28226
rect 9138 28102 9758 28170
rect 9138 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 9758 28102
rect 9138 27978 9758 28046
rect 9138 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 9758 27978
rect 9138 10350 9758 27922
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 9138 -1120 9758 9922
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 597212 36758 598268
rect 36138 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 36758 597212
rect 36138 597088 36758 597156
rect 36138 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 36758 597088
rect 36138 596964 36758 597032
rect 36138 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 36758 596964
rect 36138 596840 36758 596908
rect 36138 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 36758 596840
rect 36138 580350 36758 596784
rect 36138 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 36758 580350
rect 36138 580226 36758 580294
rect 36138 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 36758 580226
rect 36138 580102 36758 580170
rect 36138 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 36758 580102
rect 36138 579978 36758 580046
rect 36138 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 36758 579978
rect 36138 562350 36758 579922
rect 36138 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 36758 562350
rect 36138 562226 36758 562294
rect 36138 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 36758 562226
rect 36138 562102 36758 562170
rect 36138 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 36758 562102
rect 36138 561978 36758 562046
rect 36138 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 36758 561978
rect 36138 544350 36758 561922
rect 36138 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 36758 544350
rect 36138 544226 36758 544294
rect 36138 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 36758 544226
rect 36138 544102 36758 544170
rect 36138 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 36758 544102
rect 36138 543978 36758 544046
rect 36138 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 36758 543978
rect 36138 526350 36758 543922
rect 36138 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 36758 526350
rect 36138 526226 36758 526294
rect 36138 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 36758 526226
rect 36138 526102 36758 526170
rect 36138 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 36758 526102
rect 36138 525978 36758 526046
rect 36138 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 36758 525978
rect 36138 508350 36758 525922
rect 36138 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 36758 508350
rect 36138 508226 36758 508294
rect 36138 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 36758 508226
rect 36138 508102 36758 508170
rect 36138 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 36758 508102
rect 36138 507978 36758 508046
rect 36138 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 36758 507978
rect 36138 490350 36758 507922
rect 36138 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 36758 490350
rect 36138 490226 36758 490294
rect 36138 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 36758 490226
rect 36138 490102 36758 490170
rect 36138 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 36758 490102
rect 36138 489978 36758 490046
rect 36138 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 36758 489978
rect 36138 472350 36758 489922
rect 36138 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 36758 472350
rect 36138 472226 36758 472294
rect 36138 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 36758 472226
rect 36138 472102 36758 472170
rect 36138 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 36758 472102
rect 36138 471978 36758 472046
rect 36138 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 36758 471978
rect 36138 454350 36758 471922
rect 36138 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 36758 454350
rect 36138 454226 36758 454294
rect 36138 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 36758 454226
rect 36138 454102 36758 454170
rect 36138 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 36758 454102
rect 36138 453978 36758 454046
rect 36138 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 36758 453978
rect 36138 436350 36758 453922
rect 36138 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 36758 436350
rect 36138 436226 36758 436294
rect 36138 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 36758 436226
rect 36138 436102 36758 436170
rect 36138 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 36758 436102
rect 36138 435978 36758 436046
rect 36138 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 36758 435978
rect 36138 418350 36758 435922
rect 36138 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 36758 418350
rect 36138 418226 36758 418294
rect 36138 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 36758 418226
rect 36138 418102 36758 418170
rect 36138 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 36758 418102
rect 36138 417978 36758 418046
rect 36138 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 36758 417978
rect 36138 400350 36758 417922
rect 36138 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 36758 400350
rect 36138 400226 36758 400294
rect 36138 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 36758 400226
rect 36138 400102 36758 400170
rect 36138 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 36758 400102
rect 36138 399978 36758 400046
rect 36138 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 36758 399978
rect 36138 382350 36758 399922
rect 36138 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 36758 382350
rect 36138 382226 36758 382294
rect 36138 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 36758 382226
rect 36138 382102 36758 382170
rect 36138 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 36758 382102
rect 36138 381978 36758 382046
rect 36138 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 36758 381978
rect 36138 364350 36758 381922
rect 36138 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 36758 364350
rect 36138 364226 36758 364294
rect 36138 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 36758 364226
rect 36138 364102 36758 364170
rect 36138 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 36758 364102
rect 36138 363978 36758 364046
rect 36138 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 36758 363978
rect 36138 346350 36758 363922
rect 36138 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 36758 346350
rect 36138 346226 36758 346294
rect 36138 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 36758 346226
rect 36138 346102 36758 346170
rect 36138 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 36758 346102
rect 36138 345978 36758 346046
rect 36138 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 36758 345978
rect 36138 328350 36758 345922
rect 36138 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 36758 328350
rect 36138 328226 36758 328294
rect 36138 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 36758 328226
rect 36138 328102 36758 328170
rect 36138 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 36758 328102
rect 36138 327978 36758 328046
rect 36138 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 36758 327978
rect 36138 310350 36758 327922
rect 36138 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 36758 310350
rect 36138 310226 36758 310294
rect 36138 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 36758 310226
rect 36138 310102 36758 310170
rect 36138 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 36758 310102
rect 36138 309978 36758 310046
rect 36138 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 36758 309978
rect 36138 292350 36758 309922
rect 36138 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 36758 292350
rect 36138 292226 36758 292294
rect 36138 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 36758 292226
rect 36138 292102 36758 292170
rect 36138 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 36758 292102
rect 36138 291978 36758 292046
rect 36138 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 36758 291978
rect 36138 274350 36758 291922
rect 36138 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 36758 274350
rect 36138 274226 36758 274294
rect 36138 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 36758 274226
rect 36138 274102 36758 274170
rect 36138 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 36758 274102
rect 36138 273978 36758 274046
rect 36138 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 36758 273978
rect 36138 256350 36758 273922
rect 36138 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 36758 256350
rect 36138 256226 36758 256294
rect 36138 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 36758 256226
rect 36138 256102 36758 256170
rect 36138 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 36758 256102
rect 36138 255978 36758 256046
rect 36138 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 36758 255978
rect 36138 238350 36758 255922
rect 36138 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 36758 238350
rect 36138 238226 36758 238294
rect 36138 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 36758 238226
rect 36138 238102 36758 238170
rect 36138 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 36758 238102
rect 36138 237978 36758 238046
rect 36138 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 36758 237978
rect 36138 220350 36758 237922
rect 36138 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 36758 220350
rect 36138 220226 36758 220294
rect 36138 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 36758 220226
rect 36138 220102 36758 220170
rect 36138 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 36758 220102
rect 36138 219978 36758 220046
rect 36138 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 36758 219978
rect 36138 202350 36758 219922
rect 36138 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 36758 202350
rect 36138 202226 36758 202294
rect 36138 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 36758 202226
rect 36138 202102 36758 202170
rect 36138 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 36758 202102
rect 36138 201978 36758 202046
rect 36138 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 36758 201978
rect 36138 184350 36758 201922
rect 36138 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 36758 184350
rect 36138 184226 36758 184294
rect 36138 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 36758 184226
rect 36138 184102 36758 184170
rect 36138 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 36758 184102
rect 36138 183978 36758 184046
rect 36138 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 36758 183978
rect 36138 166350 36758 183922
rect 36138 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 36758 166350
rect 36138 166226 36758 166294
rect 36138 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 36758 166226
rect 36138 166102 36758 166170
rect 36138 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 36758 166102
rect 36138 165978 36758 166046
rect 36138 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 36758 165978
rect 36138 148350 36758 165922
rect 36138 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 36758 148350
rect 36138 148226 36758 148294
rect 36138 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 36758 148226
rect 36138 148102 36758 148170
rect 36138 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 36758 148102
rect 36138 147978 36758 148046
rect 36138 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 36758 147978
rect 36138 130350 36758 147922
rect 36138 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 36758 130350
rect 36138 130226 36758 130294
rect 36138 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 36758 130226
rect 36138 130102 36758 130170
rect 36138 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 36758 130102
rect 36138 129978 36758 130046
rect 36138 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 36758 129978
rect 36138 112350 36758 129922
rect 36138 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 36758 112350
rect 36138 112226 36758 112294
rect 36138 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 36758 112226
rect 36138 112102 36758 112170
rect 36138 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 36758 112102
rect 36138 111978 36758 112046
rect 36138 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 36758 111978
rect 36138 94350 36758 111922
rect 36138 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 36758 94350
rect 36138 94226 36758 94294
rect 36138 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 36758 94226
rect 36138 94102 36758 94170
rect 36138 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 36758 94102
rect 36138 93978 36758 94046
rect 36138 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 36758 93978
rect 36138 76350 36758 93922
rect 36138 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 36758 76350
rect 36138 76226 36758 76294
rect 36138 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 36758 76226
rect 36138 76102 36758 76170
rect 36138 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 36758 76102
rect 36138 75978 36758 76046
rect 36138 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 36758 75978
rect 36138 58350 36758 75922
rect 36138 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 36758 58350
rect 36138 58226 36758 58294
rect 36138 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 36758 58226
rect 36138 58102 36758 58170
rect 36138 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 36758 58102
rect 36138 57978 36758 58046
rect 36138 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 36758 57978
rect 36138 40350 36758 57922
rect 36138 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 36758 40350
rect 36138 40226 36758 40294
rect 36138 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 36758 40226
rect 36138 40102 36758 40170
rect 36138 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 36758 40102
rect 36138 39978 36758 40046
rect 36138 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 36758 39978
rect 36138 22350 36758 39922
rect 36138 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 36758 22350
rect 36138 22226 36758 22294
rect 36138 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 36758 22226
rect 36138 22102 36758 22170
rect 36138 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 36758 22102
rect 36138 21978 36758 22046
rect 36138 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 36758 21978
rect 36138 4350 36758 21922
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 66858 597212 67478 598268
rect 66858 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 67478 597212
rect 66858 597088 67478 597156
rect 66858 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 67478 597088
rect 66858 596964 67478 597032
rect 66858 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 67478 596964
rect 66858 596840 67478 596908
rect 66858 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 67478 596840
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 568350 40478 585922
rect 51996 588644 52052 588654
rect 39858 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 40478 568350
rect 39858 568226 40478 568294
rect 39858 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 40478 568226
rect 39858 568102 40478 568170
rect 39858 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 40478 568102
rect 39858 567978 40478 568046
rect 39858 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 40478 567978
rect 39858 550350 40478 567922
rect 39858 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 40478 550350
rect 39858 550226 40478 550294
rect 39858 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 40478 550226
rect 39858 550102 40478 550170
rect 39858 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 40478 550102
rect 39858 549978 40478 550046
rect 39858 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 40478 549978
rect 39858 532350 40478 549922
rect 39858 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532294 40478 532350
rect 39858 532226 40478 532294
rect 39858 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 40478 532226
rect 39858 532102 40478 532170
rect 39858 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 40478 532102
rect 39858 531978 40478 532046
rect 39858 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 40478 531978
rect 39858 514350 40478 531922
rect 39858 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 40478 514350
rect 39858 514226 40478 514294
rect 39858 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 40478 514226
rect 39858 514102 40478 514170
rect 39858 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 40478 514102
rect 39858 513978 40478 514046
rect 39858 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 40478 513978
rect 39858 496350 40478 513922
rect 39858 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 40478 496350
rect 39858 496226 40478 496294
rect 39858 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 40478 496226
rect 39858 496102 40478 496170
rect 39858 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 40478 496102
rect 39858 495978 40478 496046
rect 39858 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 40478 495978
rect 39858 478350 40478 495922
rect 39858 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 40478 478350
rect 39858 478226 40478 478294
rect 39858 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 40478 478226
rect 39858 478102 40478 478170
rect 39858 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 40478 478102
rect 39858 477978 40478 478046
rect 39858 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 40478 477978
rect 39858 460350 40478 477922
rect 39858 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 40478 460350
rect 39858 460226 40478 460294
rect 39858 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 40478 460226
rect 39858 460102 40478 460170
rect 39858 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 40478 460102
rect 39858 459978 40478 460046
rect 39858 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 40478 459978
rect 39858 442350 40478 459922
rect 39858 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 40478 442350
rect 39858 442226 40478 442294
rect 39858 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 40478 442226
rect 39858 442102 40478 442170
rect 39858 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 40478 442102
rect 39858 441978 40478 442046
rect 39858 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 40478 441978
rect 39858 424350 40478 441922
rect 39858 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 40478 424350
rect 39858 424226 40478 424294
rect 39858 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 40478 424226
rect 39858 424102 40478 424170
rect 39858 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 40478 424102
rect 39858 423978 40478 424046
rect 39858 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 40478 423978
rect 39858 406350 40478 423922
rect 39858 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 40478 406350
rect 39858 406226 40478 406294
rect 39858 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 40478 406226
rect 39858 406102 40478 406170
rect 39858 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 40478 406102
rect 39858 405978 40478 406046
rect 39858 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 40478 405978
rect 39858 388350 40478 405922
rect 39858 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 40478 388350
rect 39858 388226 40478 388294
rect 39858 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 40478 388226
rect 39858 388102 40478 388170
rect 39858 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 40478 388102
rect 39858 387978 40478 388046
rect 39858 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 40478 387978
rect 39858 370350 40478 387922
rect 39858 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 40478 370350
rect 39858 370226 40478 370294
rect 39858 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 40478 370226
rect 39858 370102 40478 370170
rect 39858 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 40478 370102
rect 39858 369978 40478 370046
rect 39858 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 40478 369978
rect 39858 352350 40478 369922
rect 39858 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 40478 352350
rect 39858 352226 40478 352294
rect 39858 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 40478 352226
rect 39858 352102 40478 352170
rect 39858 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 40478 352102
rect 39858 351978 40478 352046
rect 39858 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 40478 351978
rect 39858 334350 40478 351922
rect 39858 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 40478 334350
rect 39858 334226 40478 334294
rect 39858 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 40478 334226
rect 39858 334102 40478 334170
rect 39858 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 40478 334102
rect 39858 333978 40478 334046
rect 39858 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 40478 333978
rect 39858 316350 40478 333922
rect 39858 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 40478 316350
rect 39858 316226 40478 316294
rect 39858 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 40478 316226
rect 39858 316102 40478 316170
rect 39858 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 40478 316102
rect 39858 315978 40478 316046
rect 39858 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 40478 315978
rect 39858 298350 40478 315922
rect 50316 575428 50372 575438
rect 50316 312900 50372 575372
rect 51996 338436 52052 588588
rect 66858 580350 67478 596784
rect 66858 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 67478 580350
rect 66858 580226 67478 580294
rect 66858 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 67478 580226
rect 66858 580102 67478 580170
rect 66858 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 67478 580102
rect 66858 579978 67478 580046
rect 66858 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 67478 579978
rect 66858 562350 67478 579922
rect 66858 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 67478 562350
rect 66858 562226 67478 562294
rect 66858 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 67478 562226
rect 66858 562102 67478 562170
rect 66858 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 67478 562102
rect 66858 561978 67478 562046
rect 66858 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 67478 561978
rect 55356 551098 55412 551108
rect 53676 382788 53732 382798
rect 53564 378756 53620 378766
rect 53452 357252 53508 357262
rect 51996 338370 52052 338380
rect 53228 355908 53284 355918
rect 50316 312834 50372 312844
rect 53116 331716 53172 331726
rect 53116 300718 53172 331660
rect 53116 300652 53172 300662
rect 39858 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 40478 298350
rect 39858 298226 40478 298294
rect 39858 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 40478 298226
rect 39858 298102 40478 298170
rect 39858 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 40478 298102
rect 39858 297978 40478 298046
rect 39858 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 40478 297978
rect 39858 280350 40478 297922
rect 53228 293698 53284 355852
rect 53228 293632 53284 293642
rect 53340 354564 53396 354574
rect 53340 285418 53396 354508
rect 53452 287218 53508 357196
rect 53564 296938 53620 378700
rect 53564 296872 53620 296882
rect 53676 291718 53732 382732
rect 54348 381444 54404 381454
rect 54348 300358 54404 381388
rect 55020 361284 55076 361294
rect 54796 358596 54852 358606
rect 54684 349188 54740 349198
rect 54572 347844 54628 347854
rect 54460 319620 54516 319630
rect 54460 300804 54516 319564
rect 54460 300738 54516 300748
rect 54348 300292 54404 300302
rect 53676 291652 53732 291662
rect 54572 288478 54628 347788
rect 54572 288412 54628 288422
rect 53452 287152 53508 287162
rect 53340 285352 53396 285362
rect 54684 280756 54740 349132
rect 54796 290638 54852 358540
rect 54796 290572 54852 290582
rect 54908 351876 54964 351886
rect 54908 281092 54964 351820
rect 55020 290278 55076 361228
rect 55244 322308 55300 322318
rect 55020 290212 55076 290222
rect 55132 303492 55188 303502
rect 55132 282178 55188 303436
rect 55132 282112 55188 282122
rect 54908 281026 54964 281036
rect 54684 280690 54740 280700
rect 39858 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 40478 280350
rect 39858 280226 40478 280294
rect 39858 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 40478 280226
rect 39858 280102 40478 280170
rect 39858 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 40478 280102
rect 39858 279978 40478 280046
rect 39858 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 40478 279978
rect 39858 262350 40478 279922
rect 39858 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 40478 262350
rect 39858 262226 40478 262294
rect 39858 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 40478 262226
rect 39858 262102 40478 262170
rect 39858 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 40478 262102
rect 39858 261978 40478 262046
rect 39858 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 40478 261978
rect 39858 244350 40478 261922
rect 39858 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 40478 244350
rect 39858 244226 40478 244294
rect 39858 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 40478 244226
rect 39858 244102 40478 244170
rect 39858 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 40478 244102
rect 39858 243978 40478 244046
rect 39858 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 40478 243978
rect 39858 226350 40478 243922
rect 39858 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 40478 226350
rect 39858 226226 40478 226294
rect 39858 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 40478 226226
rect 39858 226102 40478 226170
rect 39858 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 40478 226102
rect 39858 225978 40478 226046
rect 39858 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 40478 225978
rect 39858 208350 40478 225922
rect 39858 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 40478 208350
rect 39858 208226 40478 208294
rect 39858 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 40478 208226
rect 39858 208102 40478 208170
rect 39858 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 40478 208102
rect 39858 207978 40478 208046
rect 39858 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 40478 207978
rect 39858 190350 40478 207922
rect 39858 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 40478 190350
rect 39858 190226 40478 190294
rect 39858 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 40478 190226
rect 39858 190102 40478 190170
rect 39858 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 40478 190102
rect 39858 189978 40478 190046
rect 39858 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 40478 189978
rect 39858 172350 40478 189922
rect 39858 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 40478 172350
rect 39858 172226 40478 172294
rect 39858 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 40478 172226
rect 39858 172102 40478 172170
rect 39858 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 40478 172102
rect 39858 171978 40478 172046
rect 39858 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 40478 171978
rect 39858 154350 40478 171922
rect 39858 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 40478 154350
rect 39858 154226 40478 154294
rect 39858 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 40478 154226
rect 39858 154102 40478 154170
rect 39858 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 40478 154102
rect 39858 153978 40478 154046
rect 39858 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 40478 153978
rect 39858 136350 40478 153922
rect 55244 145348 55300 322252
rect 55356 311556 55412 551042
rect 58716 547858 58772 547868
rect 56476 429940 56532 429950
rect 56364 427140 56420 427150
rect 56364 386820 56420 427084
rect 56476 389508 56532 429884
rect 56588 427258 56644 427268
rect 56588 413700 56644 427202
rect 57036 427078 57092 427088
rect 56588 413634 56644 413644
rect 56700 425098 56756 425108
rect 56700 392196 56756 425042
rect 56700 392130 56756 392140
rect 56812 423478 56868 423488
rect 56812 390852 56868 423422
rect 57036 412356 57092 427022
rect 57036 412290 57092 412300
rect 56812 390786 56868 390796
rect 56476 389442 56532 389452
rect 56364 386754 56420 386764
rect 56924 388164 56980 388174
rect 55356 311490 55412 311500
rect 56140 385476 56196 385486
rect 56028 302148 56084 302158
rect 55356 300916 55412 300926
rect 55356 261268 55412 300860
rect 56028 267988 56084 302092
rect 56140 292740 56196 385420
rect 56812 377412 56868 377422
rect 56700 373380 56756 373390
rect 56588 372036 56644 372046
rect 56476 362628 56532 362638
rect 56364 359940 56420 359950
rect 56140 292674 56196 292684
rect 56252 353220 56308 353230
rect 56252 291732 56308 353164
rect 56364 291956 56420 359884
rect 56476 292292 56532 362572
rect 56476 292226 56532 292236
rect 56588 292180 56644 371980
rect 56588 292114 56644 292124
rect 56364 291890 56420 291900
rect 56252 291666 56308 291676
rect 56700 291620 56756 373324
rect 56812 292068 56868 377356
rect 56924 297118 56980 388108
rect 58716 384748 58772 547802
rect 66858 544350 67478 561922
rect 66858 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 67478 544350
rect 66858 544226 67478 544294
rect 66858 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 67478 544226
rect 66858 544102 67478 544170
rect 66858 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 67478 544102
rect 66858 543978 67478 544046
rect 66858 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 67478 543978
rect 66858 533992 67478 543922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 568350 71198 585922
rect 70578 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 71198 568350
rect 70578 568226 71198 568294
rect 70578 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 71198 568226
rect 70578 568102 71198 568170
rect 70578 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 71198 568102
rect 70578 567978 71198 568046
rect 70578 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 71198 567978
rect 70578 550350 71198 567922
rect 97578 597212 98198 598268
rect 97578 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 98198 597212
rect 97578 597088 98198 597156
rect 97578 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 98198 597088
rect 97578 596964 98198 597032
rect 97578 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 98198 596964
rect 97578 596840 98198 596908
rect 97578 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 98198 596840
rect 97578 580350 98198 596784
rect 97578 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 98198 580350
rect 97578 580226 98198 580294
rect 97578 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 98198 580226
rect 97578 580102 98198 580170
rect 97578 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 98198 580102
rect 97578 579978 98198 580046
rect 97578 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 98198 579978
rect 97578 562350 98198 579922
rect 97578 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 98198 562350
rect 97578 562226 98198 562294
rect 97578 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 98198 562226
rect 97578 562102 98198 562170
rect 97578 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 98198 562102
rect 97578 561978 98198 562046
rect 97578 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 98198 561978
rect 97578 551392 98198 561922
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 101298 586350 101918 597744
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 101298 568350 101918 585922
rect 101298 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 101918 568350
rect 101298 568226 101918 568294
rect 101298 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 101918 568226
rect 101298 568102 101918 568170
rect 101298 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 101918 568102
rect 101298 567978 101918 568046
rect 101298 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 101918 567978
rect 101298 556192 101918 567922
rect 128298 597212 128918 598268
rect 128298 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 128918 597212
rect 128298 597088 128918 597156
rect 128298 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 128918 597088
rect 128298 596964 128918 597032
rect 128298 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 128918 596964
rect 128298 596840 128918 596908
rect 128298 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 128918 596840
rect 128298 580350 128918 596784
rect 128298 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 128918 580350
rect 128298 580226 128918 580294
rect 128298 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 128918 580226
rect 128298 580102 128918 580170
rect 128298 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 128918 580102
rect 128298 579978 128918 580046
rect 128298 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 128918 579978
rect 128298 562350 128918 579922
rect 128298 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 128918 562350
rect 128298 562226 128918 562294
rect 128298 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 128918 562226
rect 128298 562102 128918 562170
rect 128298 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 128918 562102
rect 128298 561978 128918 562046
rect 128298 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 128918 561978
rect 70578 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 71198 550350
rect 70578 550226 71198 550294
rect 70578 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 71198 550226
rect 70578 550102 71198 550170
rect 70578 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 71198 550102
rect 70578 549978 71198 550046
rect 70578 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 71198 549978
rect 70578 536872 71198 549922
rect 121996 548038 122052 548048
rect 94800 544433 95000 544446
rect 94800 544377 94810 544433
rect 94866 544377 94934 544433
rect 94990 544377 95000 544433
rect 94800 544309 95000 544377
rect 94800 544253 94810 544309
rect 94866 544253 94934 544309
rect 94990 544253 95000 544309
rect 94800 544240 95000 544253
rect 95048 544433 95496 544446
rect 95048 544377 95058 544433
rect 95114 544377 95182 544433
rect 95238 544377 95306 544433
rect 95362 544377 95430 544433
rect 95486 544377 95496 544433
rect 95048 544309 95496 544377
rect 95048 544253 95058 544309
rect 95114 544253 95182 544309
rect 95238 544253 95306 544309
rect 95362 544253 95430 544309
rect 95486 544253 95496 544309
rect 95048 544240 95496 544253
rect 95544 544433 95992 544446
rect 95544 544377 95554 544433
rect 95610 544377 95678 544433
rect 95734 544377 95802 544433
rect 95858 544377 95926 544433
rect 95982 544377 95992 544433
rect 95544 544309 95992 544377
rect 95544 544253 95554 544309
rect 95610 544253 95678 544309
rect 95734 544253 95802 544309
rect 95858 544253 95926 544309
rect 95982 544253 95992 544309
rect 95544 544240 95992 544253
rect 96040 544433 96488 544446
rect 96040 544377 96050 544433
rect 96106 544377 96174 544433
rect 96230 544377 96298 544433
rect 96354 544377 96422 544433
rect 96478 544377 96488 544433
rect 96040 544309 96488 544377
rect 96040 544253 96050 544309
rect 96106 544253 96174 544309
rect 96230 544253 96298 544309
rect 96354 544253 96422 544309
rect 96478 544253 96488 544309
rect 96040 544240 96488 544253
rect 96536 544433 96984 544446
rect 96536 544377 96546 544433
rect 96602 544377 96670 544433
rect 96726 544377 96794 544433
rect 96850 544377 96918 544433
rect 96974 544377 96984 544433
rect 96536 544309 96984 544377
rect 96536 544253 96546 544309
rect 96602 544253 96670 544309
rect 96726 544253 96794 544309
rect 96850 544253 96918 544309
rect 96974 544253 96984 544309
rect 96536 544240 96984 544253
rect 97032 544433 97480 544446
rect 97032 544377 97042 544433
rect 97098 544377 97166 544433
rect 97222 544377 97290 544433
rect 97346 544377 97414 544433
rect 97470 544377 97480 544433
rect 97032 544309 97480 544377
rect 97032 544253 97042 544309
rect 97098 544253 97166 544309
rect 97222 544253 97290 544309
rect 97346 544253 97414 544309
rect 97470 544253 97480 544309
rect 97032 544240 97480 544253
rect 97528 544433 97976 544446
rect 97528 544377 97538 544433
rect 97594 544377 97662 544433
rect 97718 544377 97786 544433
rect 97842 544377 97910 544433
rect 97966 544377 97976 544433
rect 97528 544309 97976 544377
rect 97528 544253 97538 544309
rect 97594 544253 97662 544309
rect 97718 544253 97786 544309
rect 97842 544253 97910 544309
rect 97966 544253 97976 544309
rect 97528 544240 97976 544253
rect 98024 544433 98472 544446
rect 98024 544377 98034 544433
rect 98090 544377 98158 544433
rect 98214 544377 98282 544433
rect 98338 544377 98406 544433
rect 98462 544377 98472 544433
rect 98024 544309 98472 544377
rect 98024 544253 98034 544309
rect 98090 544253 98158 544309
rect 98214 544253 98282 544309
rect 98338 544253 98406 544309
rect 98462 544253 98472 544309
rect 98024 544240 98472 544253
rect 98520 544433 98968 544446
rect 98520 544377 98530 544433
rect 98586 544377 98654 544433
rect 98710 544377 98778 544433
rect 98834 544377 98902 544433
rect 98958 544377 98968 544433
rect 98520 544309 98968 544377
rect 98520 544253 98530 544309
rect 98586 544253 98654 544309
rect 98710 544253 98778 544309
rect 98834 544253 98902 544309
rect 98958 544253 98968 544309
rect 98520 544240 98968 544253
rect 99016 544433 99464 544446
rect 99016 544377 99026 544433
rect 99082 544377 99150 544433
rect 99206 544377 99274 544433
rect 99330 544377 99398 544433
rect 99454 544377 99464 544433
rect 99016 544309 99464 544377
rect 99016 544253 99026 544309
rect 99082 544253 99150 544309
rect 99206 544253 99274 544309
rect 99330 544253 99398 544309
rect 99454 544253 99464 544309
rect 99016 544240 99464 544253
rect 99512 544433 99960 544446
rect 99512 544377 99522 544433
rect 99578 544377 99646 544433
rect 99702 544377 99770 544433
rect 99826 544377 99894 544433
rect 99950 544377 99960 544433
rect 99512 544309 99960 544377
rect 99512 544253 99522 544309
rect 99578 544253 99646 544309
rect 99702 544253 99770 544309
rect 99826 544253 99894 544309
rect 99950 544253 99960 544309
rect 99512 544240 99960 544253
rect 100008 544433 100456 544446
rect 100008 544377 100018 544433
rect 100074 544377 100142 544433
rect 100198 544377 100266 544433
rect 100322 544377 100390 544433
rect 100446 544377 100456 544433
rect 100008 544309 100456 544377
rect 100008 544253 100018 544309
rect 100074 544253 100142 544309
rect 100198 544253 100266 544309
rect 100322 544253 100390 544309
rect 100446 544253 100456 544309
rect 100008 544240 100456 544253
rect 100504 544433 100952 544446
rect 100504 544377 100514 544433
rect 100570 544377 100638 544433
rect 100694 544377 100762 544433
rect 100818 544377 100886 544433
rect 100942 544377 100952 544433
rect 100504 544309 100952 544377
rect 100504 544253 100514 544309
rect 100570 544253 100638 544309
rect 100694 544253 100762 544309
rect 100818 544253 100886 544309
rect 100942 544253 100952 544309
rect 100504 544240 100952 544253
rect 101000 544433 101448 544446
rect 101000 544377 101010 544433
rect 101066 544377 101134 544433
rect 101190 544377 101258 544433
rect 101314 544377 101382 544433
rect 101438 544377 101448 544433
rect 101000 544309 101448 544377
rect 101000 544253 101010 544309
rect 101066 544253 101134 544309
rect 101190 544253 101258 544309
rect 101314 544253 101382 544309
rect 101438 544253 101448 544309
rect 101000 544240 101448 544253
rect 101496 544433 101944 544446
rect 101496 544377 101506 544433
rect 101562 544377 101630 544433
rect 101686 544377 101754 544433
rect 101810 544377 101878 544433
rect 101934 544377 101944 544433
rect 101496 544309 101944 544377
rect 101496 544253 101506 544309
rect 101562 544253 101630 544309
rect 101686 544253 101754 544309
rect 101810 544253 101878 544309
rect 101934 544253 101944 544309
rect 101496 544240 101944 544253
rect 101992 544433 102440 544446
rect 101992 544377 102002 544433
rect 102058 544377 102126 544433
rect 102182 544377 102250 544433
rect 102306 544377 102374 544433
rect 102430 544377 102440 544433
rect 101992 544309 102440 544377
rect 101992 544253 102002 544309
rect 102058 544253 102126 544309
rect 102182 544253 102250 544309
rect 102306 544253 102374 544309
rect 102430 544253 102440 544309
rect 101992 544240 102440 544253
rect 102488 544433 102936 544446
rect 102488 544377 102498 544433
rect 102554 544377 102622 544433
rect 102678 544377 102746 544433
rect 102802 544377 102870 544433
rect 102926 544377 102936 544433
rect 102488 544309 102936 544377
rect 102488 544253 102498 544309
rect 102554 544253 102622 544309
rect 102678 544253 102746 544309
rect 102802 544253 102870 544309
rect 102926 544253 102936 544309
rect 102488 544240 102936 544253
rect 102984 544433 103432 544446
rect 102984 544377 102994 544433
rect 103050 544377 103118 544433
rect 103174 544377 103242 544433
rect 103298 544377 103366 544433
rect 103422 544377 103432 544433
rect 102984 544309 103432 544377
rect 102984 544253 102994 544309
rect 103050 544253 103118 544309
rect 103174 544253 103242 544309
rect 103298 544253 103366 544309
rect 103422 544253 103432 544309
rect 102984 544240 103432 544253
rect 103480 544433 103928 544446
rect 103480 544377 103490 544433
rect 103546 544377 103614 544433
rect 103670 544377 103738 544433
rect 103794 544377 103862 544433
rect 103918 544377 103928 544433
rect 103480 544309 103928 544377
rect 103480 544253 103490 544309
rect 103546 544253 103614 544309
rect 103670 544253 103738 544309
rect 103794 544253 103862 544309
rect 103918 544253 103928 544309
rect 103480 544240 103928 544253
rect 103976 544433 104424 544446
rect 103976 544377 103986 544433
rect 104042 544377 104110 544433
rect 104166 544377 104234 544433
rect 104290 544377 104358 544433
rect 104414 544377 104424 544433
rect 103976 544309 104424 544377
rect 103976 544253 103986 544309
rect 104042 544253 104110 544309
rect 104166 544253 104234 544309
rect 104290 544253 104358 544309
rect 104414 544253 104424 544309
rect 103976 544240 104424 544253
rect 104472 544433 104920 544446
rect 104472 544377 104482 544433
rect 104538 544377 104606 544433
rect 104662 544377 104730 544433
rect 104786 544377 104854 544433
rect 104910 544377 104920 544433
rect 104472 544309 104920 544377
rect 104472 544253 104482 544309
rect 104538 544253 104606 544309
rect 104662 544253 104730 544309
rect 104786 544253 104854 544309
rect 104910 544253 104920 544309
rect 104472 544240 104920 544253
rect 104968 544433 105416 544446
rect 104968 544377 104978 544433
rect 105034 544377 105102 544433
rect 105158 544377 105226 544433
rect 105282 544377 105350 544433
rect 105406 544377 105416 544433
rect 104968 544309 105416 544377
rect 104968 544253 104978 544309
rect 105034 544253 105102 544309
rect 105158 544253 105226 544309
rect 105282 544253 105350 544309
rect 105406 544253 105416 544309
rect 104968 544240 105416 544253
rect 105464 544433 105912 544446
rect 105464 544377 105474 544433
rect 105530 544377 105598 544433
rect 105654 544377 105722 544433
rect 105778 544377 105846 544433
rect 105902 544377 105912 544433
rect 105464 544309 105912 544377
rect 105464 544253 105474 544309
rect 105530 544253 105598 544309
rect 105654 544253 105722 544309
rect 105778 544253 105846 544309
rect 105902 544253 105912 544309
rect 105464 544240 105912 544253
rect 105960 544433 106408 544446
rect 105960 544377 105970 544433
rect 106026 544377 106094 544433
rect 106150 544377 106218 544433
rect 106274 544377 106342 544433
rect 106398 544377 106408 544433
rect 105960 544309 106408 544377
rect 105960 544253 105970 544309
rect 106026 544253 106094 544309
rect 106150 544253 106218 544309
rect 106274 544253 106342 544309
rect 106398 544253 106408 544309
rect 105960 544240 106408 544253
rect 106456 544433 106904 544446
rect 106456 544377 106466 544433
rect 106522 544377 106590 544433
rect 106646 544377 106714 544433
rect 106770 544377 106838 544433
rect 106894 544377 106904 544433
rect 106456 544309 106904 544377
rect 106456 544253 106466 544309
rect 106522 544253 106590 544309
rect 106646 544253 106714 544309
rect 106770 544253 106838 544309
rect 106894 544253 106904 544309
rect 106456 544240 106904 544253
rect 106952 544433 107400 544446
rect 106952 544377 106962 544433
rect 107018 544377 107086 544433
rect 107142 544377 107210 544433
rect 107266 544377 107334 544433
rect 107390 544377 107400 544433
rect 106952 544309 107400 544377
rect 106952 544253 106962 544309
rect 107018 544253 107086 544309
rect 107142 544253 107210 544309
rect 107266 544253 107334 544309
rect 107390 544253 107400 544309
rect 106952 544240 107400 544253
rect 94560 544090 107280 544120
rect 94560 544034 94630 544090
rect 94686 544034 94754 544090
rect 94810 544034 94878 544090
rect 94934 544034 95002 544090
rect 95058 544034 95126 544090
rect 95182 544034 95250 544090
rect 95306 544034 95374 544090
rect 95430 544034 95498 544090
rect 95554 544034 95622 544090
rect 95678 544034 95746 544090
rect 95802 544034 95870 544090
rect 95926 544034 95994 544090
rect 96050 544034 96118 544090
rect 96174 544034 96242 544090
rect 96298 544034 96366 544090
rect 96422 544034 96490 544090
rect 96546 544034 96614 544090
rect 96670 544034 96738 544090
rect 96794 544034 96862 544090
rect 96918 544034 96986 544090
rect 97042 544034 97110 544090
rect 97166 544034 97234 544090
rect 97290 544034 97358 544090
rect 97414 544034 97482 544090
rect 97538 544034 97606 544090
rect 97662 544034 97730 544090
rect 97786 544034 97854 544090
rect 97910 544034 97978 544090
rect 98034 544034 98102 544090
rect 98158 544034 98226 544090
rect 98282 544034 98350 544090
rect 98406 544034 98474 544090
rect 98530 544034 98598 544090
rect 98654 544034 98722 544090
rect 98778 544034 98846 544090
rect 98902 544034 98970 544090
rect 99026 544034 99094 544090
rect 99150 544034 99218 544090
rect 99274 544034 99342 544090
rect 99398 544034 99466 544090
rect 99522 544034 99590 544090
rect 99646 544034 99714 544090
rect 99770 544034 99838 544090
rect 99894 544034 99962 544090
rect 100018 544034 100086 544090
rect 100142 544034 100210 544090
rect 100266 544034 100334 544090
rect 100390 544034 100458 544090
rect 100514 544034 100582 544090
rect 100638 544034 100706 544090
rect 100762 544034 100830 544090
rect 100886 544034 100954 544090
rect 101010 544034 101078 544090
rect 101134 544034 101202 544090
rect 101258 544034 101326 544090
rect 101382 544034 101450 544090
rect 101506 544034 101574 544090
rect 101630 544034 101698 544090
rect 101754 544034 101822 544090
rect 101878 544034 101946 544090
rect 102002 544034 102070 544090
rect 102126 544034 102194 544090
rect 102250 544034 102318 544090
rect 102374 544034 102442 544090
rect 102498 544034 102566 544090
rect 102622 544034 102690 544090
rect 102746 544034 102814 544090
rect 102870 544034 102938 544090
rect 102994 544034 103062 544090
rect 103118 544034 103186 544090
rect 103242 544034 103310 544090
rect 103366 544034 103434 544090
rect 103490 544034 103558 544090
rect 103614 544034 103682 544090
rect 103738 544034 103806 544090
rect 103862 544034 103930 544090
rect 103986 544034 104054 544090
rect 104110 544034 104178 544090
rect 104234 544034 104302 544090
rect 104358 544034 104426 544090
rect 104482 544034 104550 544090
rect 104606 544034 104674 544090
rect 104730 544034 104798 544090
rect 104854 544034 104922 544090
rect 104978 544034 105046 544090
rect 105102 544034 105170 544090
rect 105226 544034 105294 544090
rect 105350 544034 105418 544090
rect 105474 544034 105542 544090
rect 105598 544034 105666 544090
rect 105722 544034 105790 544090
rect 105846 544034 105914 544090
rect 105970 544034 106038 544090
rect 106094 544034 106162 544090
rect 106218 544034 106286 544090
rect 106342 544034 106410 544090
rect 106466 544034 106534 544090
rect 106590 544034 106658 544090
rect 106714 544034 106782 544090
rect 106838 544034 106906 544090
rect 106962 544034 107030 544090
rect 107086 544034 107154 544090
rect 107210 544034 107280 544090
rect 94560 543966 107280 544034
rect 94560 543910 94630 543966
rect 94686 543910 94754 543966
rect 94810 543910 94878 543966
rect 94934 543910 95002 543966
rect 95058 543910 95126 543966
rect 95182 543910 95250 543966
rect 95306 543910 95374 543966
rect 95430 543910 95498 543966
rect 95554 543910 95622 543966
rect 95678 543910 95746 543966
rect 95802 543910 95870 543966
rect 95926 543910 95994 543966
rect 96050 543910 96118 543966
rect 96174 543910 96242 543966
rect 96298 543910 96366 543966
rect 96422 543910 96490 543966
rect 96546 543910 96614 543966
rect 96670 543910 96738 543966
rect 96794 543910 96862 543966
rect 96918 543910 96986 543966
rect 97042 543910 97110 543966
rect 97166 543910 97234 543966
rect 97290 543910 97358 543966
rect 97414 543910 97482 543966
rect 97538 543910 97606 543966
rect 97662 543910 97730 543966
rect 97786 543910 97854 543966
rect 97910 543910 97978 543966
rect 98034 543910 98102 543966
rect 98158 543910 98226 543966
rect 98282 543910 98350 543966
rect 98406 543910 98474 543966
rect 98530 543910 98598 543966
rect 98654 543910 98722 543966
rect 98778 543910 98846 543966
rect 98902 543910 98970 543966
rect 99026 543910 99094 543966
rect 99150 543910 99218 543966
rect 99274 543910 99342 543966
rect 99398 543910 99466 543966
rect 99522 543910 99590 543966
rect 99646 543910 99714 543966
rect 99770 543910 99838 543966
rect 99894 543910 99962 543966
rect 100018 543910 100086 543966
rect 100142 543910 100210 543966
rect 100266 543910 100334 543966
rect 100390 543910 100458 543966
rect 100514 543910 100582 543966
rect 100638 543910 100706 543966
rect 100762 543910 100830 543966
rect 100886 543910 100954 543966
rect 101010 543910 101078 543966
rect 101134 543910 101202 543966
rect 101258 543910 101326 543966
rect 101382 543910 101450 543966
rect 101506 543910 101574 543966
rect 101630 543910 101698 543966
rect 101754 543910 101822 543966
rect 101878 543910 101946 543966
rect 102002 543910 102070 543966
rect 102126 543910 102194 543966
rect 102250 543910 102318 543966
rect 102374 543910 102442 543966
rect 102498 543910 102566 543966
rect 102622 543910 102690 543966
rect 102746 543910 102814 543966
rect 102870 543910 102938 543966
rect 102994 543910 103062 543966
rect 103118 543910 103186 543966
rect 103242 543910 103310 543966
rect 103366 543910 103434 543966
rect 103490 543910 103558 543966
rect 103614 543910 103682 543966
rect 103738 543910 103806 543966
rect 103862 543910 103930 543966
rect 103986 543910 104054 543966
rect 104110 543910 104178 543966
rect 104234 543910 104302 543966
rect 104358 543910 104426 543966
rect 104482 543910 104550 543966
rect 104606 543910 104674 543966
rect 104730 543910 104798 543966
rect 104854 543910 104922 543966
rect 104978 543910 105046 543966
rect 105102 543910 105170 543966
rect 105226 543910 105294 543966
rect 105350 543910 105418 543966
rect 105474 543910 105542 543966
rect 105598 543910 105666 543966
rect 105722 543910 105790 543966
rect 105846 543910 105914 543966
rect 105970 543910 106038 543966
rect 106094 543910 106162 543966
rect 106218 543910 106286 543966
rect 106342 543910 106410 543966
rect 106466 543910 106534 543966
rect 106590 543910 106658 543966
rect 106714 543910 106782 543966
rect 106838 543910 106906 543966
rect 106962 543910 107030 543966
rect 107086 543910 107154 543966
rect 107210 543910 107280 543966
rect 94560 543880 107280 543910
rect 68040 532328 75480 532360
rect 68040 532272 68074 532328
rect 68130 532272 68198 532328
rect 68254 532272 68322 532328
rect 68378 532272 68446 532328
rect 68502 532272 68570 532328
rect 68626 532272 68694 532328
rect 68750 532272 68818 532328
rect 68874 532272 68942 532328
rect 68998 532272 69066 532328
rect 69122 532272 69190 532328
rect 69246 532272 69314 532328
rect 69370 532272 69438 532328
rect 69494 532272 69562 532328
rect 69618 532272 69686 532328
rect 69742 532272 69810 532328
rect 69866 532272 69934 532328
rect 69990 532272 70058 532328
rect 70114 532272 70182 532328
rect 70238 532272 70306 532328
rect 70362 532272 70430 532328
rect 70486 532272 70554 532328
rect 70610 532272 70678 532328
rect 70734 532272 70802 532328
rect 70858 532272 70926 532328
rect 70982 532272 71050 532328
rect 71106 532272 71174 532328
rect 71230 532272 71298 532328
rect 71354 532272 71422 532328
rect 71478 532272 71546 532328
rect 71602 532272 71670 532328
rect 71726 532272 71794 532328
rect 71850 532272 71918 532328
rect 71974 532272 72042 532328
rect 72098 532272 72166 532328
rect 72222 532272 72290 532328
rect 72346 532272 72414 532328
rect 72470 532272 72538 532328
rect 72594 532272 72662 532328
rect 72718 532272 72786 532328
rect 72842 532272 72910 532328
rect 72966 532272 73034 532328
rect 73090 532272 73158 532328
rect 73214 532272 73282 532328
rect 73338 532272 73406 532328
rect 73462 532272 73530 532328
rect 73586 532272 73654 532328
rect 73710 532272 73778 532328
rect 73834 532272 73902 532328
rect 73958 532272 74026 532328
rect 74082 532272 74150 532328
rect 74206 532272 74274 532328
rect 74330 532272 74398 532328
rect 74454 532272 74522 532328
rect 74578 532272 74646 532328
rect 74702 532272 74770 532328
rect 74826 532272 74894 532328
rect 74950 532272 75018 532328
rect 75074 532272 75142 532328
rect 75198 532272 75266 532328
rect 75322 532272 75390 532328
rect 75446 532272 75480 532328
rect 68040 532240 75480 532272
rect 84840 526328 98760 526360
rect 84840 526272 84890 526328
rect 84946 526272 85014 526328
rect 85070 526272 85138 526328
rect 85194 526272 85262 526328
rect 85318 526272 85386 526328
rect 85442 526272 85510 526328
rect 85566 526272 85634 526328
rect 85690 526272 85758 526328
rect 85814 526272 85882 526328
rect 85938 526272 86006 526328
rect 86062 526272 86130 526328
rect 86186 526272 86254 526328
rect 86310 526272 86378 526328
rect 86434 526272 86502 526328
rect 86558 526272 86626 526328
rect 86682 526272 86750 526328
rect 86806 526272 86874 526328
rect 86930 526272 86998 526328
rect 87054 526272 87122 526328
rect 87178 526272 87246 526328
rect 87302 526272 87370 526328
rect 87426 526272 87494 526328
rect 87550 526272 87618 526328
rect 87674 526272 87742 526328
rect 87798 526272 87866 526328
rect 87922 526272 87990 526328
rect 88046 526272 88114 526328
rect 88170 526272 88238 526328
rect 88294 526272 88362 526328
rect 88418 526272 88486 526328
rect 88542 526272 88610 526328
rect 88666 526272 88734 526328
rect 88790 526272 88858 526328
rect 88914 526272 88982 526328
rect 89038 526272 89106 526328
rect 89162 526272 89230 526328
rect 89286 526272 89354 526328
rect 89410 526272 89478 526328
rect 89534 526272 89602 526328
rect 89658 526272 89726 526328
rect 89782 526272 89850 526328
rect 89906 526272 89974 526328
rect 90030 526272 90098 526328
rect 90154 526272 90222 526328
rect 90278 526272 90346 526328
rect 90402 526272 90470 526328
rect 90526 526272 90594 526328
rect 90650 526272 90718 526328
rect 90774 526272 90842 526328
rect 90898 526272 90966 526328
rect 91022 526272 91090 526328
rect 91146 526272 91214 526328
rect 91270 526272 91338 526328
rect 91394 526272 91462 526328
rect 91518 526272 91586 526328
rect 91642 526272 91710 526328
rect 91766 526272 91834 526328
rect 91890 526272 91958 526328
rect 92014 526272 92082 526328
rect 92138 526272 92206 526328
rect 92262 526272 92330 526328
rect 92386 526272 92454 526328
rect 92510 526272 92578 526328
rect 92634 526272 92702 526328
rect 92758 526272 92826 526328
rect 92882 526272 92950 526328
rect 93006 526272 93074 526328
rect 93130 526272 93198 526328
rect 93254 526272 93322 526328
rect 93378 526272 93446 526328
rect 93502 526272 93570 526328
rect 93626 526272 93694 526328
rect 93750 526272 93818 526328
rect 93874 526272 93942 526328
rect 93998 526272 94066 526328
rect 94122 526272 94190 526328
rect 94246 526272 94314 526328
rect 94370 526272 94438 526328
rect 94494 526272 94562 526328
rect 94618 526272 94686 526328
rect 94742 526272 94810 526328
rect 94866 526272 94934 526328
rect 94990 526272 95058 526328
rect 95114 526272 95182 526328
rect 95238 526272 95306 526328
rect 95362 526272 95430 526328
rect 95486 526272 95554 526328
rect 95610 526272 95678 526328
rect 95734 526272 95802 526328
rect 95858 526272 95926 526328
rect 95982 526272 96050 526328
rect 96106 526272 96174 526328
rect 96230 526272 96298 526328
rect 96354 526272 96422 526328
rect 96478 526272 96546 526328
rect 96602 526272 96670 526328
rect 96726 526272 96794 526328
rect 96850 526272 96918 526328
rect 96974 526272 97042 526328
rect 97098 526272 97166 526328
rect 97222 526272 97290 526328
rect 97346 526272 97414 526328
rect 97470 526272 97538 526328
rect 97594 526272 97662 526328
rect 97718 526272 97786 526328
rect 97842 526272 97910 526328
rect 97966 526272 98034 526328
rect 98090 526272 98158 526328
rect 98214 526272 98282 526328
rect 98338 526272 98406 526328
rect 98462 526272 98530 526328
rect 98586 526272 98654 526328
rect 98710 526272 98760 526328
rect 84840 526240 98760 526272
rect 84720 526090 98520 526120
rect 84720 526034 84772 526090
rect 84828 526034 84896 526090
rect 84952 526034 85020 526090
rect 85076 526034 85144 526090
rect 85200 526034 85268 526090
rect 85324 526034 85392 526090
rect 85448 526034 85516 526090
rect 85572 526034 85640 526090
rect 85696 526034 85764 526090
rect 85820 526034 85888 526090
rect 85944 526034 86012 526090
rect 86068 526034 86136 526090
rect 86192 526034 86260 526090
rect 86316 526034 86384 526090
rect 86440 526034 86508 526090
rect 86564 526034 86632 526090
rect 86688 526034 86756 526090
rect 86812 526034 86880 526090
rect 86936 526034 87004 526090
rect 87060 526034 87128 526090
rect 87184 526034 87252 526090
rect 87308 526034 87376 526090
rect 87432 526034 87500 526090
rect 87556 526034 87624 526090
rect 87680 526034 87748 526090
rect 87804 526034 87872 526090
rect 87928 526034 87996 526090
rect 88052 526034 88120 526090
rect 88176 526034 88244 526090
rect 88300 526034 88368 526090
rect 88424 526034 88492 526090
rect 88548 526034 88616 526090
rect 88672 526034 88740 526090
rect 88796 526034 88864 526090
rect 88920 526034 88988 526090
rect 89044 526034 89112 526090
rect 89168 526034 89236 526090
rect 89292 526034 89360 526090
rect 89416 526034 89484 526090
rect 89540 526034 89608 526090
rect 89664 526034 89732 526090
rect 89788 526034 89856 526090
rect 89912 526034 89980 526090
rect 90036 526034 90104 526090
rect 90160 526034 90228 526090
rect 90284 526034 90352 526090
rect 90408 526034 90476 526090
rect 90532 526034 90600 526090
rect 90656 526034 90724 526090
rect 90780 526034 90848 526090
rect 90904 526034 90972 526090
rect 91028 526034 91096 526090
rect 91152 526034 91220 526090
rect 91276 526034 91344 526090
rect 91400 526034 91468 526090
rect 91524 526034 91592 526090
rect 91648 526034 91716 526090
rect 91772 526034 91840 526090
rect 91896 526034 91964 526090
rect 92020 526034 92088 526090
rect 92144 526034 92212 526090
rect 92268 526034 92336 526090
rect 92392 526034 92460 526090
rect 92516 526034 92584 526090
rect 92640 526034 92708 526090
rect 92764 526034 92832 526090
rect 92888 526034 92956 526090
rect 93012 526034 93080 526090
rect 93136 526034 93204 526090
rect 93260 526034 93328 526090
rect 93384 526034 93452 526090
rect 93508 526034 93576 526090
rect 93632 526034 93700 526090
rect 93756 526034 93824 526090
rect 93880 526034 93948 526090
rect 94004 526034 94072 526090
rect 94128 526034 94196 526090
rect 94252 526034 94320 526090
rect 94376 526034 94444 526090
rect 94500 526034 94568 526090
rect 94624 526034 94692 526090
rect 94748 526034 94816 526090
rect 94872 526034 94940 526090
rect 94996 526034 95064 526090
rect 95120 526034 95188 526090
rect 95244 526034 95312 526090
rect 95368 526034 95436 526090
rect 95492 526034 95560 526090
rect 95616 526034 95684 526090
rect 95740 526034 95808 526090
rect 95864 526034 95932 526090
rect 95988 526034 96056 526090
rect 96112 526034 96180 526090
rect 96236 526034 96304 526090
rect 96360 526034 96428 526090
rect 96484 526034 96552 526090
rect 96608 526034 96676 526090
rect 96732 526034 96800 526090
rect 96856 526034 96924 526090
rect 96980 526034 97048 526090
rect 97104 526034 97172 526090
rect 97228 526034 97296 526090
rect 97352 526034 97420 526090
rect 97476 526034 97544 526090
rect 97600 526034 97668 526090
rect 97724 526034 97792 526090
rect 97848 526034 97916 526090
rect 97972 526034 98040 526090
rect 98096 526034 98164 526090
rect 98220 526034 98288 526090
rect 98344 526034 98412 526090
rect 98468 526034 98520 526090
rect 84720 525966 98520 526034
rect 84720 525910 84772 525966
rect 84828 525910 84896 525966
rect 84952 525910 85020 525966
rect 85076 525910 85144 525966
rect 85200 525910 85268 525966
rect 85324 525910 85392 525966
rect 85448 525910 85516 525966
rect 85572 525910 85640 525966
rect 85696 525910 85764 525966
rect 85820 525910 85888 525966
rect 85944 525910 86012 525966
rect 86068 525910 86136 525966
rect 86192 525910 86260 525966
rect 86316 525910 86384 525966
rect 86440 525910 86508 525966
rect 86564 525910 86632 525966
rect 86688 525910 86756 525966
rect 86812 525910 86880 525966
rect 86936 525910 87004 525966
rect 87060 525910 87128 525966
rect 87184 525910 87252 525966
rect 87308 525910 87376 525966
rect 87432 525910 87500 525966
rect 87556 525910 87624 525966
rect 87680 525910 87748 525966
rect 87804 525910 87872 525966
rect 87928 525910 87996 525966
rect 88052 525910 88120 525966
rect 88176 525910 88244 525966
rect 88300 525910 88368 525966
rect 88424 525910 88492 525966
rect 88548 525910 88616 525966
rect 88672 525910 88740 525966
rect 88796 525910 88864 525966
rect 88920 525910 88988 525966
rect 89044 525910 89112 525966
rect 89168 525910 89236 525966
rect 89292 525910 89360 525966
rect 89416 525910 89484 525966
rect 89540 525910 89608 525966
rect 89664 525910 89732 525966
rect 89788 525910 89856 525966
rect 89912 525910 89980 525966
rect 90036 525910 90104 525966
rect 90160 525910 90228 525966
rect 90284 525910 90352 525966
rect 90408 525910 90476 525966
rect 90532 525910 90600 525966
rect 90656 525910 90724 525966
rect 90780 525910 90848 525966
rect 90904 525910 90972 525966
rect 91028 525910 91096 525966
rect 91152 525910 91220 525966
rect 91276 525910 91344 525966
rect 91400 525910 91468 525966
rect 91524 525910 91592 525966
rect 91648 525910 91716 525966
rect 91772 525910 91840 525966
rect 91896 525910 91964 525966
rect 92020 525910 92088 525966
rect 92144 525910 92212 525966
rect 92268 525910 92336 525966
rect 92392 525910 92460 525966
rect 92516 525910 92584 525966
rect 92640 525910 92708 525966
rect 92764 525910 92832 525966
rect 92888 525910 92956 525966
rect 93012 525910 93080 525966
rect 93136 525910 93204 525966
rect 93260 525910 93328 525966
rect 93384 525910 93452 525966
rect 93508 525910 93576 525966
rect 93632 525910 93700 525966
rect 93756 525910 93824 525966
rect 93880 525910 93948 525966
rect 94004 525910 94072 525966
rect 94128 525910 94196 525966
rect 94252 525910 94320 525966
rect 94376 525910 94444 525966
rect 94500 525910 94568 525966
rect 94624 525910 94692 525966
rect 94748 525910 94816 525966
rect 94872 525910 94940 525966
rect 94996 525910 95064 525966
rect 95120 525910 95188 525966
rect 95244 525910 95312 525966
rect 95368 525910 95436 525966
rect 95492 525910 95560 525966
rect 95616 525910 95684 525966
rect 95740 525910 95808 525966
rect 95864 525910 95932 525966
rect 95988 525910 96056 525966
rect 96112 525910 96180 525966
rect 96236 525910 96304 525966
rect 96360 525910 96428 525966
rect 96484 525910 96552 525966
rect 96608 525910 96676 525966
rect 96732 525910 96800 525966
rect 96856 525910 96924 525966
rect 96980 525910 97048 525966
rect 97104 525910 97172 525966
rect 97228 525910 97296 525966
rect 97352 525910 97420 525966
rect 97476 525910 97544 525966
rect 97600 525910 97668 525966
rect 97724 525910 97792 525966
rect 97848 525910 97916 525966
rect 97972 525910 98040 525966
rect 98096 525910 98164 525966
rect 98220 525910 98288 525966
rect 98344 525910 98412 525966
rect 98468 525910 98520 525966
rect 84720 525880 98520 525910
rect 60000 514412 60232 514446
rect 60000 514356 60026 514412
rect 60082 514356 60150 514412
rect 60206 514356 60232 514412
rect 60000 514288 60232 514356
rect 60000 514232 60026 514288
rect 60082 514232 60150 514288
rect 60206 514232 60232 514288
rect 60000 514164 60232 514232
rect 60000 514108 60026 514164
rect 60082 514108 60150 514164
rect 60206 514108 60232 514164
rect 60000 514040 60232 514108
rect 60000 513984 60026 514040
rect 60082 513984 60150 514040
rect 60206 513984 60232 514040
rect 60000 513916 60232 513984
rect 60000 513860 60026 513916
rect 60082 513860 60150 513916
rect 60206 513860 60232 513916
rect 60000 513826 60232 513860
rect 60248 514412 60728 514446
rect 60248 514356 60274 514412
rect 60330 514356 60398 514412
rect 60454 514356 60522 514412
rect 60578 514356 60646 514412
rect 60702 514356 60728 514412
rect 60248 514288 60728 514356
rect 60248 514232 60274 514288
rect 60330 514232 60398 514288
rect 60454 514232 60522 514288
rect 60578 514232 60646 514288
rect 60702 514232 60728 514288
rect 60248 514164 60728 514232
rect 60248 514108 60274 514164
rect 60330 514108 60398 514164
rect 60454 514108 60522 514164
rect 60578 514108 60646 514164
rect 60702 514108 60728 514164
rect 60248 514040 60728 514108
rect 60248 513984 60274 514040
rect 60330 513984 60398 514040
rect 60454 513984 60522 514040
rect 60578 513984 60646 514040
rect 60702 513984 60728 514040
rect 60248 513916 60728 513984
rect 60248 513860 60274 513916
rect 60330 513860 60398 513916
rect 60454 513860 60522 513916
rect 60578 513860 60646 513916
rect 60702 513860 60728 513916
rect 60248 513826 60728 513860
rect 60744 514412 61224 514446
rect 60744 514356 60770 514412
rect 60826 514356 60894 514412
rect 60950 514356 61018 514412
rect 61074 514356 61142 514412
rect 61198 514356 61224 514412
rect 60744 514288 61224 514356
rect 60744 514232 60770 514288
rect 60826 514232 60894 514288
rect 60950 514232 61018 514288
rect 61074 514232 61142 514288
rect 61198 514232 61224 514288
rect 60744 514164 61224 514232
rect 60744 514108 60770 514164
rect 60826 514108 60894 514164
rect 60950 514108 61018 514164
rect 61074 514108 61142 514164
rect 61198 514108 61224 514164
rect 60744 514040 61224 514108
rect 60744 513984 60770 514040
rect 60826 513984 60894 514040
rect 60950 513984 61018 514040
rect 61074 513984 61142 514040
rect 61198 513984 61224 514040
rect 60744 513916 61224 513984
rect 60744 513860 60770 513916
rect 60826 513860 60894 513916
rect 60950 513860 61018 513916
rect 61074 513860 61142 513916
rect 61198 513860 61224 513916
rect 60744 513826 61224 513860
rect 61240 514412 61720 514446
rect 61240 514356 61266 514412
rect 61322 514356 61390 514412
rect 61446 514356 61514 514412
rect 61570 514356 61638 514412
rect 61694 514356 61720 514412
rect 61240 514288 61720 514356
rect 61240 514232 61266 514288
rect 61322 514232 61390 514288
rect 61446 514232 61514 514288
rect 61570 514232 61638 514288
rect 61694 514232 61720 514288
rect 61240 514164 61720 514232
rect 61240 514108 61266 514164
rect 61322 514108 61390 514164
rect 61446 514108 61514 514164
rect 61570 514108 61638 514164
rect 61694 514108 61720 514164
rect 61240 514040 61720 514108
rect 61240 513984 61266 514040
rect 61322 513984 61390 514040
rect 61446 513984 61514 514040
rect 61570 513984 61638 514040
rect 61694 513984 61720 514040
rect 61240 513916 61720 513984
rect 61240 513860 61266 513916
rect 61322 513860 61390 513916
rect 61446 513860 61514 513916
rect 61570 513860 61638 513916
rect 61694 513860 61720 513916
rect 61240 513826 61720 513860
rect 61736 514412 62216 514446
rect 61736 514356 61762 514412
rect 61818 514356 61886 514412
rect 61942 514356 62010 514412
rect 62066 514356 62134 514412
rect 62190 514356 62216 514412
rect 61736 514288 62216 514356
rect 61736 514232 61762 514288
rect 61818 514232 61886 514288
rect 61942 514232 62010 514288
rect 62066 514232 62134 514288
rect 62190 514232 62216 514288
rect 61736 514164 62216 514232
rect 61736 514108 61762 514164
rect 61818 514108 61886 514164
rect 61942 514108 62010 514164
rect 62066 514108 62134 514164
rect 62190 514108 62216 514164
rect 61736 514040 62216 514108
rect 61736 513984 61762 514040
rect 61818 513984 61886 514040
rect 61942 513984 62010 514040
rect 62066 513984 62134 514040
rect 62190 513984 62216 514040
rect 61736 513916 62216 513984
rect 61736 513860 61762 513916
rect 61818 513860 61886 513916
rect 61942 513860 62010 513916
rect 62066 513860 62134 513916
rect 62190 513860 62216 513916
rect 61736 513826 62216 513860
rect 62232 514412 62712 514446
rect 62232 514356 62258 514412
rect 62314 514356 62382 514412
rect 62438 514356 62506 514412
rect 62562 514356 62630 514412
rect 62686 514356 62712 514412
rect 62232 514288 62712 514356
rect 62232 514232 62258 514288
rect 62314 514232 62382 514288
rect 62438 514232 62506 514288
rect 62562 514232 62630 514288
rect 62686 514232 62712 514288
rect 62232 514164 62712 514232
rect 62232 514108 62258 514164
rect 62314 514108 62382 514164
rect 62438 514108 62506 514164
rect 62562 514108 62630 514164
rect 62686 514108 62712 514164
rect 62232 514040 62712 514108
rect 62232 513984 62258 514040
rect 62314 513984 62382 514040
rect 62438 513984 62506 514040
rect 62562 513984 62630 514040
rect 62686 513984 62712 514040
rect 62232 513916 62712 513984
rect 62232 513860 62258 513916
rect 62314 513860 62382 513916
rect 62438 513860 62506 513916
rect 62562 513860 62630 513916
rect 62686 513860 62712 513916
rect 62232 513826 62712 513860
rect 62728 514412 63208 514446
rect 62728 514356 62754 514412
rect 62810 514356 62878 514412
rect 62934 514356 63002 514412
rect 63058 514356 63126 514412
rect 63182 514356 63208 514412
rect 62728 514288 63208 514356
rect 62728 514232 62754 514288
rect 62810 514232 62878 514288
rect 62934 514232 63002 514288
rect 63058 514232 63126 514288
rect 63182 514232 63208 514288
rect 62728 514164 63208 514232
rect 62728 514108 62754 514164
rect 62810 514108 62878 514164
rect 62934 514108 63002 514164
rect 63058 514108 63126 514164
rect 63182 514108 63208 514164
rect 62728 514040 63208 514108
rect 62728 513984 62754 514040
rect 62810 513984 62878 514040
rect 62934 513984 63002 514040
rect 63058 513984 63126 514040
rect 63182 513984 63208 514040
rect 62728 513916 63208 513984
rect 62728 513860 62754 513916
rect 62810 513860 62878 513916
rect 62934 513860 63002 513916
rect 63058 513860 63126 513916
rect 63182 513860 63208 513916
rect 62728 513826 63208 513860
rect 63224 514412 63704 514446
rect 63224 514356 63250 514412
rect 63306 514356 63374 514412
rect 63430 514356 63498 514412
rect 63554 514356 63622 514412
rect 63678 514356 63704 514412
rect 63224 514288 63704 514356
rect 63224 514232 63250 514288
rect 63306 514232 63374 514288
rect 63430 514232 63498 514288
rect 63554 514232 63622 514288
rect 63678 514232 63704 514288
rect 63224 514164 63704 514232
rect 63224 514108 63250 514164
rect 63306 514108 63374 514164
rect 63430 514108 63498 514164
rect 63554 514108 63622 514164
rect 63678 514108 63704 514164
rect 63224 514040 63704 514108
rect 63224 513984 63250 514040
rect 63306 513984 63374 514040
rect 63430 513984 63498 514040
rect 63554 513984 63622 514040
rect 63678 513984 63704 514040
rect 63224 513916 63704 513984
rect 63224 513860 63250 513916
rect 63306 513860 63374 513916
rect 63430 513860 63498 513916
rect 63554 513860 63622 513916
rect 63678 513860 63704 513916
rect 63224 513826 63704 513860
rect 63720 514412 64200 514446
rect 63720 514356 63746 514412
rect 63802 514356 63870 514412
rect 63926 514356 63994 514412
rect 64050 514356 64118 514412
rect 64174 514356 64200 514412
rect 63720 514288 64200 514356
rect 63720 514232 63746 514288
rect 63802 514232 63870 514288
rect 63926 514232 63994 514288
rect 64050 514232 64118 514288
rect 64174 514232 64200 514288
rect 63720 514164 64200 514232
rect 63720 514108 63746 514164
rect 63802 514108 63870 514164
rect 63926 514108 63994 514164
rect 64050 514108 64118 514164
rect 64174 514108 64200 514164
rect 63720 514040 64200 514108
rect 63720 513984 63746 514040
rect 63802 513984 63870 514040
rect 63926 513984 63994 514040
rect 64050 513984 64118 514040
rect 64174 513984 64200 514040
rect 63720 513916 64200 513984
rect 63720 513860 63746 513916
rect 63802 513860 63870 513916
rect 63926 513860 63994 513916
rect 64050 513860 64118 513916
rect 64174 513860 64200 513916
rect 63720 513826 64200 513860
rect 78960 508431 79160 508446
rect 78960 508375 78970 508431
rect 79026 508375 79094 508431
rect 79150 508375 79160 508431
rect 78960 508360 79160 508375
rect 79208 508431 79656 508446
rect 79208 508375 79218 508431
rect 79274 508375 79342 508431
rect 79398 508375 79466 508431
rect 79522 508375 79590 508431
rect 79646 508375 79656 508431
rect 79208 508360 79656 508375
rect 79704 508431 80152 508446
rect 79704 508375 79714 508431
rect 79770 508375 79838 508431
rect 79894 508375 79962 508431
rect 80018 508375 80086 508431
rect 80142 508375 80152 508431
rect 79704 508360 80152 508375
rect 80200 508431 80648 508446
rect 80200 508375 80210 508431
rect 80266 508375 80334 508431
rect 80390 508375 80458 508431
rect 80514 508375 80582 508431
rect 80638 508375 80648 508431
rect 80200 508360 80648 508375
rect 80696 508431 81144 508446
rect 80696 508375 80706 508431
rect 80762 508375 80830 508431
rect 80886 508375 80954 508431
rect 81010 508375 81078 508431
rect 81134 508375 81144 508431
rect 80696 508360 81144 508375
rect 81192 508431 81640 508446
rect 81192 508375 81202 508431
rect 81258 508375 81326 508431
rect 81382 508375 81450 508431
rect 81506 508375 81574 508431
rect 81630 508375 81640 508431
rect 81192 508360 81640 508375
rect 81688 508431 82136 508446
rect 81688 508375 81698 508431
rect 81754 508375 81822 508431
rect 81878 508375 81946 508431
rect 82002 508375 82070 508431
rect 82126 508375 82136 508431
rect 81688 508360 82136 508375
rect 82184 508431 82632 508446
rect 82184 508375 82194 508431
rect 82250 508375 82318 508431
rect 82374 508375 82442 508431
rect 82498 508375 82566 508431
rect 82622 508375 82632 508431
rect 82184 508360 82632 508375
rect 82680 508431 83128 508446
rect 82680 508375 82690 508431
rect 82746 508375 82814 508431
rect 82870 508375 82938 508431
rect 82994 508375 83062 508431
rect 83118 508375 83128 508431
rect 82680 508360 83128 508375
rect 83176 508431 83624 508446
rect 83176 508375 83186 508431
rect 83242 508375 83310 508431
rect 83366 508375 83434 508431
rect 83490 508375 83558 508431
rect 83614 508375 83624 508431
rect 83176 508360 83624 508375
rect 83672 508431 84120 508446
rect 83672 508375 83682 508431
rect 83738 508375 83806 508431
rect 83862 508375 83930 508431
rect 83986 508375 84054 508431
rect 84110 508375 84120 508431
rect 83672 508360 84120 508375
rect 78840 508208 79040 508240
rect 78840 508152 78850 508208
rect 78906 508152 78974 508208
rect 79030 508152 79040 508208
rect 78840 508120 79040 508152
rect 79088 508208 79536 508240
rect 79088 508152 79098 508208
rect 79154 508152 79222 508208
rect 79278 508152 79346 508208
rect 79402 508152 79470 508208
rect 79526 508152 79536 508208
rect 79088 508120 79536 508152
rect 79584 508208 80032 508240
rect 79584 508152 79594 508208
rect 79650 508152 79718 508208
rect 79774 508152 79842 508208
rect 79898 508152 79966 508208
rect 80022 508152 80032 508208
rect 79584 508120 80032 508152
rect 80080 508208 80528 508240
rect 80080 508152 80090 508208
rect 80146 508152 80214 508208
rect 80270 508152 80338 508208
rect 80394 508152 80462 508208
rect 80518 508152 80528 508208
rect 80080 508120 80528 508152
rect 80576 508208 81024 508240
rect 80576 508152 80586 508208
rect 80642 508152 80710 508208
rect 80766 508152 80834 508208
rect 80890 508152 80958 508208
rect 81014 508152 81024 508208
rect 80576 508120 81024 508152
rect 81072 508208 81520 508240
rect 81072 508152 81082 508208
rect 81138 508152 81206 508208
rect 81262 508152 81330 508208
rect 81386 508152 81454 508208
rect 81510 508152 81520 508208
rect 81072 508120 81520 508152
rect 81568 508208 82016 508240
rect 81568 508152 81578 508208
rect 81634 508152 81702 508208
rect 81758 508152 81826 508208
rect 81882 508152 81950 508208
rect 82006 508152 82016 508208
rect 81568 508120 82016 508152
rect 82064 508208 82512 508240
rect 82064 508152 82074 508208
rect 82130 508152 82198 508208
rect 82254 508152 82322 508208
rect 82378 508152 82446 508208
rect 82502 508152 82512 508208
rect 82064 508120 82512 508152
rect 82560 508208 83008 508240
rect 82560 508152 82570 508208
rect 82626 508152 82694 508208
rect 82750 508152 82818 508208
rect 82874 508152 82942 508208
rect 82998 508152 83008 508208
rect 82560 508120 83008 508152
rect 83056 508208 83504 508240
rect 83056 508152 83066 508208
rect 83122 508152 83190 508208
rect 83246 508152 83314 508208
rect 83370 508152 83438 508208
rect 83494 508152 83504 508208
rect 83056 508120 83504 508152
rect 83552 508208 84000 508240
rect 83552 508152 83562 508208
rect 83618 508152 83686 508208
rect 83742 508152 83810 508208
rect 83866 508152 83934 508208
rect 83990 508152 84000 508208
rect 83552 508120 84000 508152
rect 67920 496328 74760 496360
rect 67920 496272 67964 496328
rect 68020 496272 68088 496328
rect 68144 496272 68212 496328
rect 68268 496272 68336 496328
rect 68392 496272 68460 496328
rect 68516 496272 68584 496328
rect 68640 496272 68708 496328
rect 68764 496272 68832 496328
rect 68888 496272 68956 496328
rect 69012 496272 69080 496328
rect 69136 496272 69204 496328
rect 69260 496272 69328 496328
rect 69384 496272 69452 496328
rect 69508 496272 69576 496328
rect 69632 496272 69700 496328
rect 69756 496272 69824 496328
rect 69880 496272 69948 496328
rect 70004 496272 70072 496328
rect 70128 496272 70196 496328
rect 70252 496272 70320 496328
rect 70376 496272 70444 496328
rect 70500 496272 70568 496328
rect 70624 496272 70692 496328
rect 70748 496272 70816 496328
rect 70872 496272 70940 496328
rect 70996 496272 71064 496328
rect 71120 496272 71188 496328
rect 71244 496272 71312 496328
rect 71368 496272 71436 496328
rect 71492 496272 71560 496328
rect 71616 496272 71684 496328
rect 71740 496272 71808 496328
rect 71864 496272 71932 496328
rect 71988 496272 72056 496328
rect 72112 496272 72180 496328
rect 72236 496272 72304 496328
rect 72360 496272 72428 496328
rect 72484 496272 72552 496328
rect 72608 496272 72676 496328
rect 72732 496272 72800 496328
rect 72856 496272 72924 496328
rect 72980 496272 73048 496328
rect 73104 496272 73172 496328
rect 73228 496272 73296 496328
rect 73352 496272 73420 496328
rect 73476 496272 73544 496328
rect 73600 496272 73668 496328
rect 73724 496272 73792 496328
rect 73848 496272 73916 496328
rect 73972 496272 74040 496328
rect 74096 496272 74164 496328
rect 74220 496272 74288 496328
rect 74344 496272 74412 496328
rect 74468 496272 74536 496328
rect 74592 496272 74660 496328
rect 74716 496272 74760 496328
rect 67920 496240 74760 496272
rect 68160 496088 74760 496120
rect 68160 496032 68208 496088
rect 68264 496032 68332 496088
rect 68388 496032 68456 496088
rect 68512 496032 68580 496088
rect 68636 496032 68704 496088
rect 68760 496032 68828 496088
rect 68884 496032 68952 496088
rect 69008 496032 69076 496088
rect 69132 496032 69200 496088
rect 69256 496032 69324 496088
rect 69380 496032 69448 496088
rect 69504 496032 69572 496088
rect 69628 496032 69696 496088
rect 69752 496032 69820 496088
rect 69876 496032 69944 496088
rect 70000 496032 70068 496088
rect 70124 496032 70192 496088
rect 70248 496032 70316 496088
rect 70372 496032 70440 496088
rect 70496 496032 70564 496088
rect 70620 496032 70688 496088
rect 70744 496032 70812 496088
rect 70868 496032 70936 496088
rect 70992 496032 71060 496088
rect 71116 496032 71184 496088
rect 71240 496032 71308 496088
rect 71364 496032 71432 496088
rect 71488 496032 71556 496088
rect 71612 496032 71680 496088
rect 71736 496032 71804 496088
rect 71860 496032 71928 496088
rect 71984 496032 72052 496088
rect 72108 496032 72176 496088
rect 72232 496032 72300 496088
rect 72356 496032 72424 496088
rect 72480 496032 72548 496088
rect 72604 496032 72672 496088
rect 72728 496032 72796 496088
rect 72852 496032 72920 496088
rect 72976 496032 73044 496088
rect 73100 496032 73168 496088
rect 73224 496032 73292 496088
rect 73348 496032 73416 496088
rect 73472 496032 73540 496088
rect 73596 496032 73664 496088
rect 73720 496032 73788 496088
rect 73844 496032 73912 496088
rect 73968 496032 74036 496088
rect 74092 496032 74160 496088
rect 74216 496032 74284 496088
rect 74340 496032 74408 496088
rect 74464 496032 74532 496088
rect 74588 496032 74656 496088
rect 74712 496032 74760 496088
rect 68160 496000 74760 496032
rect 66858 490350 67478 494488
rect 66858 490294 66954 490350
rect 67010 490294 67078 490350
rect 67134 490294 67202 490350
rect 67258 490294 67326 490350
rect 67382 490294 67478 490350
rect 66858 490226 67478 490294
rect 66858 490170 66954 490226
rect 67010 490170 67078 490226
rect 67134 490170 67202 490226
rect 67258 490170 67326 490226
rect 67382 490170 67478 490226
rect 66858 490102 67478 490170
rect 66858 490046 66954 490102
rect 67010 490046 67078 490102
rect 67134 490046 67202 490102
rect 67258 490046 67326 490102
rect 67382 490046 67478 490102
rect 66858 489978 67478 490046
rect 66858 489922 66954 489978
rect 67010 489922 67078 489978
rect 67134 489922 67202 489978
rect 67258 489922 67326 489978
rect 67382 489922 67478 489978
rect 63756 476308 63812 476318
rect 60620 428596 60676 428606
rect 60172 409798 60228 409808
rect 60172 409220 60228 409742
rect 60172 409154 60228 409164
rect 60284 408178 60340 408188
rect 60284 407764 60340 408122
rect 60284 407698 60340 407708
rect 60508 404758 60564 404768
rect 60508 404664 60564 404684
rect 58604 384692 58772 384748
rect 57932 380100 57988 380110
rect 57036 306180 57092 306190
rect 57036 300804 57092 306124
rect 57932 301798 57988 380044
rect 58604 372988 58660 384692
rect 60284 383348 60340 383358
rect 60284 383158 60340 383292
rect 60284 383092 60340 383102
rect 60172 375396 60228 375406
rect 60172 374698 60228 375340
rect 60172 374632 60228 374642
rect 58604 372932 58772 372988
rect 58492 365316 58548 365326
rect 58156 329028 58212 329038
rect 57932 301732 57988 301742
rect 58044 323652 58100 323662
rect 57036 300738 57092 300748
rect 56924 297052 56980 297062
rect 56812 292002 56868 292012
rect 56924 295428 56980 295438
rect 56700 291554 56756 291564
rect 56924 271348 56980 295372
rect 56924 271282 56980 271292
rect 56028 267922 56084 267932
rect 55356 261202 55412 261212
rect 58044 152516 58100 323596
rect 58156 295678 58212 328972
rect 58156 295612 58212 295622
rect 58268 326340 58324 326350
rect 58268 278068 58324 326284
rect 58268 278002 58324 278012
rect 58380 320964 58436 320974
rect 58380 273028 58436 320908
rect 58492 296758 58548 365260
rect 58716 337092 58772 372932
rect 60172 368676 60228 368686
rect 60172 368218 60228 368620
rect 60172 368152 60228 368162
rect 58716 337026 58772 337036
rect 60060 363972 60116 363982
rect 58716 310212 58772 310222
rect 58492 296692 58548 296702
rect 58604 308868 58660 308878
rect 58604 281998 58660 308812
rect 58716 295498 58772 310156
rect 58716 295432 58772 295442
rect 60060 283618 60116 363916
rect 60508 350084 60564 350094
rect 60508 349972 60564 349982
rect 60284 346500 60340 346510
rect 60172 335998 60228 336008
rect 60172 335076 60228 335942
rect 60172 335010 60228 335020
rect 60172 329476 60228 329486
rect 60172 329338 60228 329420
rect 60172 329272 60228 329282
rect 60284 314188 60340 346444
rect 60508 344484 60564 344496
rect 60508 344392 60564 344402
rect 60508 333060 60564 333070
rect 60396 324324 60452 324336
rect 60396 324232 60452 324242
rect 60172 314132 60340 314188
rect 60172 287038 60228 314132
rect 60284 304836 60340 304846
rect 60284 288838 60340 304780
rect 60508 301618 60564 333004
rect 60508 301552 60564 301562
rect 60284 288772 60340 288782
rect 60508 296772 60564 296782
rect 60172 286972 60228 286982
rect 60060 283552 60116 283562
rect 58604 281932 58660 281942
rect 58380 272962 58436 272972
rect 60508 160580 60564 296716
rect 60620 278292 60676 428540
rect 60732 374878 60788 374888
rect 60732 374724 60788 374822
rect 60732 374658 60788 374668
rect 60732 368038 60788 368048
rect 60732 367938 60788 367948
rect 60732 366660 60788 366670
rect 60732 366418 60788 366604
rect 60732 366352 60788 366362
rect 60732 335818 60788 335828
rect 60732 335748 60788 335762
rect 60732 335682 60788 335692
rect 60732 327684 60788 327694
rect 60732 326818 60788 327628
rect 60732 326752 60788 326762
rect 60732 307558 60788 307568
rect 60732 307458 60788 307468
rect 63756 290164 63812 476252
rect 66858 472350 67478 489922
rect 66858 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 67478 472350
rect 66858 472226 67478 472294
rect 66858 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 67478 472226
rect 66858 472102 67478 472170
rect 66858 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 67478 472102
rect 66858 471978 67478 472046
rect 66858 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 67478 471978
rect 66858 454350 67478 471922
rect 66858 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 67478 454350
rect 66858 454226 67478 454294
rect 66858 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 67478 454226
rect 66858 454102 67478 454170
rect 66858 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 67478 454102
rect 66858 453978 67478 454046
rect 66858 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 67478 453978
rect 66858 436350 67478 453922
rect 66858 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 67478 436350
rect 66858 436226 67478 436294
rect 66858 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 67478 436226
rect 66858 436102 67478 436170
rect 66858 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 67478 436102
rect 66858 435978 67478 436046
rect 66858 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 67478 435978
rect 66668 430052 66724 430062
rect 64448 418350 64768 418384
rect 64448 418294 64518 418350
rect 64574 418294 64642 418350
rect 64698 418294 64768 418350
rect 64448 418226 64768 418294
rect 64448 418170 64518 418226
rect 64574 418170 64642 418226
rect 64698 418170 64768 418226
rect 64448 418102 64768 418170
rect 64448 418046 64518 418102
rect 64574 418046 64642 418102
rect 64698 418046 64768 418102
rect 64448 417978 64768 418046
rect 64448 417922 64518 417978
rect 64574 417922 64642 417978
rect 64698 417922 64768 417978
rect 64448 417888 64768 417922
rect 64448 400350 64768 400384
rect 64448 400294 64518 400350
rect 64574 400294 64642 400350
rect 64698 400294 64768 400350
rect 64448 400226 64768 400294
rect 64448 400170 64518 400226
rect 64574 400170 64642 400226
rect 64698 400170 64768 400226
rect 64448 400102 64768 400170
rect 64448 400046 64518 400102
rect 64574 400046 64642 400102
rect 64698 400046 64768 400102
rect 64448 399978 64768 400046
rect 64448 399922 64518 399978
rect 64574 399922 64642 399978
rect 64698 399922 64768 399978
rect 64448 399888 64768 399922
rect 64448 382350 64768 382384
rect 64448 382294 64518 382350
rect 64574 382294 64642 382350
rect 64698 382294 64768 382350
rect 64448 382226 64768 382294
rect 64448 382170 64518 382226
rect 64574 382170 64642 382226
rect 64698 382170 64768 382226
rect 64448 382102 64768 382170
rect 64448 382046 64518 382102
rect 64574 382046 64642 382102
rect 64698 382046 64768 382102
rect 64448 381978 64768 382046
rect 64448 381922 64518 381978
rect 64574 381922 64642 381978
rect 64698 381922 64768 381978
rect 64448 381888 64768 381922
rect 64448 364350 64768 364384
rect 64448 364294 64518 364350
rect 64574 364294 64642 364350
rect 64698 364294 64768 364350
rect 64448 364226 64768 364294
rect 64448 364170 64518 364226
rect 64574 364170 64642 364226
rect 64698 364170 64768 364226
rect 64448 364102 64768 364170
rect 64448 364046 64518 364102
rect 64574 364046 64642 364102
rect 64698 364046 64768 364102
rect 64448 363978 64768 364046
rect 64448 363922 64518 363978
rect 64574 363922 64642 363978
rect 64698 363922 64768 363978
rect 64448 363888 64768 363922
rect 64448 346350 64768 346384
rect 64448 346294 64518 346350
rect 64574 346294 64642 346350
rect 64698 346294 64768 346350
rect 64448 346226 64768 346294
rect 64448 346170 64518 346226
rect 64574 346170 64642 346226
rect 64698 346170 64768 346226
rect 64448 346102 64768 346170
rect 64448 346046 64518 346102
rect 64574 346046 64642 346102
rect 64698 346046 64768 346102
rect 64448 345978 64768 346046
rect 64448 345922 64518 345978
rect 64574 345922 64642 345978
rect 64698 345922 64768 345978
rect 64448 345888 64768 345922
rect 64448 328350 64768 328384
rect 64448 328294 64518 328350
rect 64574 328294 64642 328350
rect 64698 328294 64768 328350
rect 64448 328226 64768 328294
rect 64448 328170 64518 328226
rect 64574 328170 64642 328226
rect 64698 328170 64768 328226
rect 64448 328102 64768 328170
rect 64448 328046 64518 328102
rect 64574 328046 64642 328102
rect 64698 328046 64768 328102
rect 64448 327978 64768 328046
rect 64448 327922 64518 327978
rect 64574 327922 64642 327978
rect 64698 327922 64768 327978
rect 64448 327888 64768 327922
rect 64448 310350 64768 310384
rect 64448 310294 64518 310350
rect 64574 310294 64642 310350
rect 64698 310294 64768 310350
rect 64448 310226 64768 310294
rect 64448 310170 64518 310226
rect 64574 310170 64642 310226
rect 64698 310170 64768 310226
rect 64448 310102 64768 310170
rect 64448 310046 64518 310102
rect 64574 310046 64642 310102
rect 64698 310046 64768 310102
rect 64448 309978 64768 310046
rect 64448 309922 64518 309978
rect 64574 309922 64642 309978
rect 64698 309922 64768 309978
rect 64448 309888 64768 309922
rect 63756 290098 63812 290108
rect 60620 278226 60676 278236
rect 66668 213332 66724 429996
rect 66668 213266 66724 213276
rect 66858 418350 67478 435922
rect 70578 478350 71198 491608
rect 70578 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 71198 478350
rect 70578 478226 71198 478294
rect 70578 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 71198 478226
rect 70578 478102 71198 478170
rect 70578 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 71198 478102
rect 70578 477978 71198 478046
rect 70578 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 71198 477978
rect 70578 460350 71198 477922
rect 70578 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 71198 460350
rect 70578 460226 71198 460294
rect 70578 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 71198 460226
rect 70578 460102 71198 460170
rect 70578 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 71198 460102
rect 70578 459978 71198 460046
rect 70578 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 71198 459978
rect 70578 442350 71198 459922
rect 70578 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 71198 442350
rect 70578 442226 71198 442294
rect 70578 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 71198 442226
rect 70578 442102 71198 442170
rect 70578 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 71198 442102
rect 70578 441978 71198 442046
rect 70578 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 71198 441978
rect 69468 431038 69524 431048
rect 69468 430276 69524 430982
rect 69468 430210 69524 430220
rect 66858 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 67478 418350
rect 66858 418226 67478 418294
rect 66858 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 67478 418226
rect 66858 418102 67478 418170
rect 66858 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 67478 418102
rect 66858 417978 67478 418046
rect 66858 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 67478 417978
rect 66858 400350 67478 417922
rect 66858 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 67478 400350
rect 66858 400226 67478 400294
rect 66858 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 67478 400226
rect 66858 400102 67478 400170
rect 66858 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 67478 400102
rect 66858 399978 67478 400046
rect 66858 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 67478 399978
rect 66858 382350 67478 399922
rect 66858 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 67478 382350
rect 66858 382226 67478 382294
rect 66858 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 67478 382226
rect 66858 382102 67478 382170
rect 66858 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 67478 382102
rect 66858 381978 67478 382046
rect 66858 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 67478 381978
rect 66858 364350 67478 381922
rect 66858 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 67478 364350
rect 66858 364226 67478 364294
rect 66858 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 67478 364226
rect 66858 364102 67478 364170
rect 66858 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 67478 364102
rect 66858 363978 67478 364046
rect 66858 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 67478 363978
rect 66858 346350 67478 363922
rect 70578 424350 71198 441922
rect 97578 490350 98198 490648
rect 97578 490294 97674 490350
rect 97730 490294 97798 490350
rect 97854 490294 97922 490350
rect 97978 490294 98046 490350
rect 98102 490294 98198 490350
rect 97578 490226 98198 490294
rect 97578 490170 97674 490226
rect 97730 490170 97798 490226
rect 97854 490170 97922 490226
rect 97978 490170 98046 490226
rect 98102 490170 98198 490226
rect 97578 490102 98198 490170
rect 97578 490046 97674 490102
rect 97730 490046 97798 490102
rect 97854 490046 97922 490102
rect 97978 490046 98046 490102
rect 98102 490046 98198 490102
rect 97578 489978 98198 490046
rect 97578 489922 97674 489978
rect 97730 489922 97798 489978
rect 97854 489922 97922 489978
rect 97978 489922 98046 489978
rect 98102 489922 98198 489978
rect 97578 472350 98198 489922
rect 97578 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 98198 472350
rect 97578 472226 98198 472294
rect 97578 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 98198 472226
rect 97578 472102 98198 472170
rect 97578 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 98198 472102
rect 97578 471978 98198 472046
rect 97578 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 98198 471978
rect 97578 454350 98198 471922
rect 97578 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 98198 454350
rect 97578 454226 98198 454294
rect 97578 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 98198 454226
rect 97578 454102 98198 454170
rect 97578 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 98198 454102
rect 97578 453978 98198 454046
rect 97578 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 98198 453978
rect 97578 436350 98198 453922
rect 97578 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 98198 436350
rect 97578 436226 98198 436294
rect 97578 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 98198 436226
rect 97578 436102 98198 436170
rect 97578 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 98198 436102
rect 97578 435978 98198 436046
rect 97578 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 98198 435978
rect 82908 432118 82964 432128
rect 76412 432068 76468 432078
rect 74844 429418 74900 429428
rect 74844 429314 74900 429324
rect 70578 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 71198 424350
rect 70578 424226 71198 424294
rect 70578 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 71198 424226
rect 70578 424102 71198 424170
rect 70578 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 71198 424102
rect 70578 423978 71198 424046
rect 70578 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 71198 423978
rect 70578 406350 71198 423922
rect 70578 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 71198 406350
rect 70578 406226 71198 406294
rect 70578 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 71198 406226
rect 70578 406102 71198 406170
rect 70578 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 71198 406102
rect 70578 405978 71198 406046
rect 70578 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 71198 405978
rect 70578 388350 71198 405922
rect 70578 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 71198 388350
rect 70578 388226 71198 388294
rect 70578 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 71198 388226
rect 70578 388102 71198 388170
rect 70578 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 71198 388102
rect 70578 387978 71198 388046
rect 70578 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 71198 387978
rect 70578 370350 71198 387922
rect 70578 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 71198 370350
rect 70578 370226 71198 370294
rect 70578 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 71198 370226
rect 70578 370102 71198 370170
rect 70578 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 71198 370102
rect 70578 369978 71198 370046
rect 70578 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 71198 369978
rect 70578 352350 71198 369922
rect 70578 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 71198 352350
rect 70578 352226 71198 352294
rect 70578 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 71198 352226
rect 70578 352102 71198 352170
rect 70578 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 71198 352102
rect 70578 351978 71198 352046
rect 70578 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 71198 351978
rect 66858 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 67478 346350
rect 66858 346226 67478 346294
rect 66858 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 67478 346226
rect 66858 346102 67478 346170
rect 66858 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 67478 346102
rect 66858 345978 67478 346046
rect 66858 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 67478 345978
rect 66858 328350 67478 345922
rect 66858 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 67478 328350
rect 66858 328226 67478 328294
rect 66858 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 67478 328226
rect 66858 328102 67478 328170
rect 66858 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 67478 328102
rect 66858 327978 67478 328046
rect 66858 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 67478 327978
rect 66858 310350 67478 327922
rect 66858 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 67478 310350
rect 66858 310226 67478 310294
rect 66858 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 67478 310226
rect 66858 310102 67478 310170
rect 66858 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 67478 310102
rect 66858 309978 67478 310046
rect 66858 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 67478 309978
rect 66858 292350 67478 309922
rect 66858 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 67478 292350
rect 66858 292226 67478 292294
rect 66858 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 67478 292226
rect 66858 292102 67478 292170
rect 66858 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 67478 292102
rect 66858 291978 67478 292046
rect 66858 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 67478 291978
rect 66858 274350 67478 291922
rect 69692 350038 69748 350048
rect 69692 290458 69748 349982
rect 69692 290392 69748 290402
rect 70578 334350 71198 351922
rect 70578 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 71198 334350
rect 70578 334226 71198 334294
rect 70578 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 71198 334226
rect 70578 334102 71198 334170
rect 70578 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 71198 334102
rect 70578 333978 71198 334046
rect 70578 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 71198 333978
rect 70578 316350 71198 333922
rect 74732 326818 74788 326828
rect 70578 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 71198 316350
rect 70578 316226 71198 316294
rect 70578 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 71198 316226
rect 70578 316102 71198 316170
rect 70578 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 71198 316102
rect 70578 315978 71198 316046
rect 70578 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 71198 315978
rect 70578 298350 71198 315922
rect 70578 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 71198 298350
rect 70578 298226 71198 298294
rect 70578 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 71198 298226
rect 70578 298102 71198 298170
rect 70578 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 71198 298102
rect 70578 297978 71198 298046
rect 70578 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 71198 297978
rect 66858 274294 66954 274350
rect 67010 274294 67078 274350
rect 67134 274294 67202 274350
rect 67258 274294 67326 274350
rect 67382 274294 67478 274350
rect 66858 274226 67478 274294
rect 66858 274170 66954 274226
rect 67010 274170 67078 274226
rect 67134 274170 67202 274226
rect 67258 274170 67326 274226
rect 67382 274170 67478 274226
rect 66858 274102 67478 274170
rect 66858 274046 66954 274102
rect 67010 274046 67078 274102
rect 67134 274046 67202 274102
rect 67258 274046 67326 274102
rect 67382 274046 67478 274102
rect 66858 273978 67478 274046
rect 66858 273922 66954 273978
rect 67010 273922 67078 273978
rect 67134 273922 67202 273978
rect 67258 273922 67326 273978
rect 67382 273922 67478 273978
rect 66858 256350 67478 273922
rect 66858 256294 66954 256350
rect 67010 256294 67078 256350
rect 67134 256294 67202 256350
rect 67258 256294 67326 256350
rect 67382 256294 67478 256350
rect 66858 256226 67478 256294
rect 66858 256170 66954 256226
rect 67010 256170 67078 256226
rect 67134 256170 67202 256226
rect 67258 256170 67326 256226
rect 67382 256170 67478 256226
rect 66858 256102 67478 256170
rect 66858 256046 66954 256102
rect 67010 256046 67078 256102
rect 67134 256046 67202 256102
rect 67258 256046 67326 256102
rect 67382 256046 67478 256102
rect 66858 255978 67478 256046
rect 66858 255922 66954 255978
rect 67010 255922 67078 255978
rect 67134 255922 67202 255978
rect 67258 255922 67326 255978
rect 67382 255922 67478 255978
rect 66858 238350 67478 255922
rect 66858 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 67478 238350
rect 66858 238226 67478 238294
rect 66858 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 67478 238226
rect 66858 238102 67478 238170
rect 66858 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 67478 238102
rect 66858 237978 67478 238046
rect 66858 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 67478 237978
rect 66858 220350 67478 237922
rect 70578 280350 71198 297922
rect 70578 280294 70674 280350
rect 70730 280294 70798 280350
rect 70854 280294 70922 280350
rect 70978 280294 71046 280350
rect 71102 280294 71198 280350
rect 70578 280226 71198 280294
rect 70578 280170 70674 280226
rect 70730 280170 70798 280226
rect 70854 280170 70922 280226
rect 70978 280170 71046 280226
rect 71102 280170 71198 280226
rect 70578 280102 71198 280170
rect 70578 280046 70674 280102
rect 70730 280046 70798 280102
rect 70854 280046 70922 280102
rect 70978 280046 71046 280102
rect 71102 280046 71198 280102
rect 70578 279978 71198 280046
rect 70578 279922 70674 279978
rect 70730 279922 70798 279978
rect 70854 279922 70922 279978
rect 70978 279922 71046 279978
rect 71102 279922 71198 279978
rect 70578 262350 71198 279922
rect 70578 262294 70674 262350
rect 70730 262294 70798 262350
rect 70854 262294 70922 262350
rect 70978 262294 71046 262350
rect 71102 262294 71198 262350
rect 70578 262226 71198 262294
rect 70578 262170 70674 262226
rect 70730 262170 70798 262226
rect 70854 262170 70922 262226
rect 70978 262170 71046 262226
rect 71102 262170 71198 262226
rect 70578 262102 71198 262170
rect 70578 262046 70674 262102
rect 70730 262046 70798 262102
rect 70854 262046 70922 262102
rect 70978 262046 71046 262102
rect 71102 262046 71198 262102
rect 70578 261978 71198 262046
rect 70578 261922 70674 261978
rect 70730 261922 70798 261978
rect 70854 261922 70922 261978
rect 70978 261922 71046 261978
rect 71102 261922 71198 261978
rect 70578 244350 71198 261922
rect 73052 324298 73108 324308
rect 73052 259588 73108 324242
rect 74732 271460 74788 326762
rect 74732 271394 74788 271404
rect 76412 264628 76468 432012
rect 82908 431956 82964 432062
rect 77532 431938 77588 431948
rect 82908 431890 82964 431900
rect 77532 431844 77588 431882
rect 77532 431778 77588 431788
rect 80220 428518 80276 428528
rect 79808 424350 80128 424384
rect 79808 424294 79878 424350
rect 79934 424294 80002 424350
rect 80058 424294 80128 424350
rect 79808 424226 80128 424294
rect 79808 424170 79878 424226
rect 79934 424170 80002 424226
rect 80058 424170 80128 424226
rect 79808 424102 80128 424170
rect 79808 424046 79878 424102
rect 79934 424046 80002 424102
rect 80058 424046 80128 424102
rect 79808 423978 80128 424046
rect 79808 423922 79878 423978
rect 79934 423922 80002 423978
rect 80058 423922 80128 423978
rect 79808 423888 80128 423922
rect 79808 406350 80128 406384
rect 79808 406294 79878 406350
rect 79934 406294 80002 406350
rect 80058 406294 80128 406350
rect 79808 406226 80128 406294
rect 79808 406170 79878 406226
rect 79934 406170 80002 406226
rect 80058 406170 80128 406226
rect 79808 406102 80128 406170
rect 79808 406046 79878 406102
rect 79934 406046 80002 406102
rect 80058 406046 80128 406102
rect 79808 405978 80128 406046
rect 79808 405922 79878 405978
rect 79934 405922 80002 405978
rect 80058 405922 80128 405978
rect 79808 405888 80128 405922
rect 79808 388350 80128 388384
rect 79808 388294 79878 388350
rect 79934 388294 80002 388350
rect 80058 388294 80128 388350
rect 79808 388226 80128 388294
rect 79808 388170 79878 388226
rect 79934 388170 80002 388226
rect 80058 388170 80128 388226
rect 79808 388102 80128 388170
rect 79808 388046 79878 388102
rect 79934 388046 80002 388102
rect 80058 388046 80128 388102
rect 79808 387978 80128 388046
rect 79808 387922 79878 387978
rect 79934 387922 80002 387978
rect 80058 387922 80128 387978
rect 79808 387888 80128 387922
rect 79808 370350 80128 370384
rect 79808 370294 79878 370350
rect 79934 370294 80002 370350
rect 80058 370294 80128 370350
rect 79808 370226 80128 370294
rect 79808 370170 79878 370226
rect 79934 370170 80002 370226
rect 80058 370170 80128 370226
rect 79808 370102 80128 370170
rect 79808 370046 79878 370102
rect 79934 370046 80002 370102
rect 80058 370046 80128 370102
rect 79808 369978 80128 370046
rect 79808 369922 79878 369978
rect 79934 369922 80002 369978
rect 80058 369922 80128 369978
rect 79808 369888 80128 369922
rect 79808 352350 80128 352384
rect 79808 352294 79878 352350
rect 79934 352294 80002 352350
rect 80058 352294 80128 352350
rect 79808 352226 80128 352294
rect 79808 352170 79878 352226
rect 79934 352170 80002 352226
rect 80058 352170 80128 352226
rect 79808 352102 80128 352170
rect 79808 352046 79878 352102
rect 79934 352046 80002 352102
rect 80058 352046 80128 352102
rect 79808 351978 80128 352046
rect 79808 351922 79878 351978
rect 79934 351922 80002 351978
rect 80058 351922 80128 351978
rect 79808 351888 80128 351922
rect 78092 344458 78148 344468
rect 76524 307558 76580 307568
rect 76524 285598 76580 307502
rect 78092 286858 78148 344402
rect 80220 335818 80276 428462
rect 83244 428484 83300 428494
rect 83132 425458 83188 425468
rect 83132 404758 83188 425402
rect 83132 404692 83188 404702
rect 80220 335752 80276 335762
rect 83132 374878 83188 374888
rect 79808 334350 80128 334384
rect 79808 334294 79878 334350
rect 79934 334294 80002 334350
rect 80058 334294 80128 334350
rect 79808 334226 80128 334294
rect 79808 334170 79878 334226
rect 79934 334170 80002 334226
rect 80058 334170 80128 334226
rect 79808 334102 80128 334170
rect 79808 334046 79878 334102
rect 79934 334046 80002 334102
rect 80058 334046 80128 334102
rect 79808 333978 80128 334046
rect 79808 333922 79878 333978
rect 79934 333922 80002 333978
rect 80058 333922 80128 333978
rect 79808 333888 80128 333922
rect 79808 316350 80128 316384
rect 79808 316294 79878 316350
rect 79934 316294 80002 316350
rect 80058 316294 80128 316350
rect 79808 316226 80128 316294
rect 79808 316170 79878 316226
rect 79934 316170 80002 316226
rect 80058 316170 80128 316226
rect 79808 316102 80128 316170
rect 79808 316046 79878 316102
rect 79934 316046 80002 316102
rect 80058 316046 80128 316102
rect 79808 315978 80128 316046
rect 79808 315922 79878 315978
rect 79934 315922 80002 315978
rect 80058 315922 80128 315978
rect 79808 315888 80128 315922
rect 79808 298350 80128 298384
rect 79808 298294 79878 298350
rect 79934 298294 80002 298350
rect 80058 298294 80128 298350
rect 79808 298226 80128 298294
rect 79808 298170 79878 298226
rect 79934 298170 80002 298226
rect 80058 298170 80128 298226
rect 79808 298102 80128 298170
rect 79808 298046 79878 298102
rect 79934 298046 80002 298102
rect 80058 298046 80128 298102
rect 79808 297978 80128 298046
rect 79808 297922 79878 297978
rect 79934 297922 80002 297978
rect 80058 297922 80128 297978
rect 79808 297888 80128 297922
rect 78092 286792 78148 286802
rect 76524 285532 76580 285542
rect 76412 264562 76468 264572
rect 81452 281428 81508 281438
rect 73052 259522 73108 259532
rect 70578 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 71198 244350
rect 70578 244226 71198 244294
rect 70578 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 71198 244226
rect 70578 244102 71198 244170
rect 70578 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 71198 244102
rect 70578 243978 71198 244046
rect 70578 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 71198 243978
rect 66858 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 67478 220350
rect 66858 220226 67478 220294
rect 66858 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 67478 220226
rect 66858 220102 67478 220170
rect 66858 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 67478 220102
rect 66858 219978 67478 220046
rect 66858 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 67478 219978
rect 62972 209972 63028 209982
rect 62972 196588 63028 209916
rect 64448 202350 64768 202384
rect 64448 202294 64518 202350
rect 64574 202294 64642 202350
rect 64698 202294 64768 202350
rect 64448 202226 64768 202294
rect 64448 202170 64518 202226
rect 64574 202170 64642 202226
rect 64698 202170 64768 202226
rect 64448 202102 64768 202170
rect 64448 202046 64518 202102
rect 64574 202046 64642 202102
rect 64698 202046 64768 202102
rect 64448 201978 64768 202046
rect 64448 201922 64518 201978
rect 64574 201922 64642 201978
rect 64698 201922 64768 201978
rect 64448 201888 64768 201922
rect 66858 202350 67478 219922
rect 66858 202294 66954 202350
rect 67010 202294 67078 202350
rect 67134 202294 67202 202350
rect 67258 202294 67326 202350
rect 67382 202294 67478 202350
rect 66858 202226 67478 202294
rect 66858 202170 66954 202226
rect 67010 202170 67078 202226
rect 67134 202170 67202 202226
rect 67258 202170 67326 202226
rect 67382 202170 67478 202226
rect 66858 202102 67478 202170
rect 66858 202046 66954 202102
rect 67010 202046 67078 202102
rect 67134 202046 67202 202102
rect 67258 202046 67326 202102
rect 67382 202046 67478 202102
rect 66858 201978 67478 202046
rect 66858 201922 66954 201978
rect 67010 201922 67078 201978
rect 67134 201922 67202 201978
rect 67258 201922 67326 201978
rect 67382 201922 67478 201978
rect 60508 160514 60564 160524
rect 62748 196532 63028 196588
rect 58044 152450 58100 152460
rect 55244 145282 55300 145292
rect 62188 142678 62244 142688
rect 62188 141988 62244 142622
rect 62748 142678 62804 196532
rect 64448 184350 64768 184384
rect 64448 184294 64518 184350
rect 64574 184294 64642 184350
rect 64698 184294 64768 184350
rect 64448 184226 64768 184294
rect 64448 184170 64518 184226
rect 64574 184170 64642 184226
rect 64698 184170 64768 184226
rect 64448 184102 64768 184170
rect 64448 184046 64518 184102
rect 64574 184046 64642 184102
rect 64698 184046 64768 184102
rect 64448 183978 64768 184046
rect 64448 183922 64518 183978
rect 64574 183922 64642 183978
rect 64698 183922 64768 183978
rect 64448 183888 64768 183922
rect 66858 184350 67478 201922
rect 66858 184294 66954 184350
rect 67010 184294 67078 184350
rect 67134 184294 67202 184350
rect 67258 184294 67326 184350
rect 67382 184294 67478 184350
rect 66858 184226 67478 184294
rect 66858 184170 66954 184226
rect 67010 184170 67078 184226
rect 67134 184170 67202 184226
rect 67258 184170 67326 184226
rect 67382 184170 67478 184226
rect 66858 184102 67478 184170
rect 66858 184046 66954 184102
rect 67010 184046 67078 184102
rect 67134 184046 67202 184102
rect 67258 184046 67326 184102
rect 67382 184046 67478 184102
rect 66858 183978 67478 184046
rect 66858 183922 66954 183978
rect 67010 183922 67078 183978
rect 67134 183922 67202 183978
rect 67258 183922 67326 183978
rect 67382 183922 67478 183978
rect 64448 166350 64768 166384
rect 64448 166294 64518 166350
rect 64574 166294 64642 166350
rect 64698 166294 64768 166350
rect 64448 166226 64768 166294
rect 64448 166170 64518 166226
rect 64574 166170 64642 166226
rect 64698 166170 64768 166226
rect 64448 166102 64768 166170
rect 64448 166046 64518 166102
rect 64574 166046 64642 166102
rect 64698 166046 64768 166102
rect 64448 165978 64768 166046
rect 64448 165922 64518 165978
rect 64574 165922 64642 165978
rect 64698 165922 64768 165978
rect 64448 165888 64768 165922
rect 66858 166350 67478 183922
rect 66858 166294 66954 166350
rect 67010 166294 67078 166350
rect 67134 166294 67202 166350
rect 67258 166294 67326 166350
rect 67382 166294 67478 166350
rect 66858 166226 67478 166294
rect 66858 166170 66954 166226
rect 67010 166170 67078 166226
rect 67134 166170 67202 166226
rect 67258 166170 67326 166226
rect 67382 166170 67478 166226
rect 66858 166102 67478 166170
rect 66858 166046 66954 166102
rect 67010 166046 67078 166102
rect 67134 166046 67202 166102
rect 67258 166046 67326 166102
rect 67382 166046 67478 166102
rect 66858 165978 67478 166046
rect 66858 165922 66954 165978
rect 67010 165922 67078 165978
rect 67134 165922 67202 165978
rect 67258 165922 67326 165978
rect 67382 165922 67478 165978
rect 62748 142612 62804 142622
rect 66858 148350 67478 165922
rect 66858 148294 66954 148350
rect 67010 148294 67078 148350
rect 67134 148294 67202 148350
rect 67258 148294 67326 148350
rect 67382 148294 67478 148350
rect 66858 148226 67478 148294
rect 66858 148170 66954 148226
rect 67010 148170 67078 148226
rect 67134 148170 67202 148226
rect 67258 148170 67326 148226
rect 67382 148170 67478 148226
rect 66858 148102 67478 148170
rect 66858 148046 66954 148102
rect 67010 148046 67078 148102
rect 67134 148046 67202 148102
rect 67258 148046 67326 148102
rect 67382 148046 67478 148102
rect 66858 147978 67478 148046
rect 66858 147922 66954 147978
rect 67010 147922 67078 147978
rect 67134 147922 67202 147978
rect 67258 147922 67326 147978
rect 67382 147922 67478 147978
rect 62188 141922 62244 141932
rect 63756 142318 63812 142328
rect 63756 141204 63812 142262
rect 63756 141138 63812 141148
rect 39858 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 40478 136350
rect 39858 136226 40478 136294
rect 39858 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 40478 136226
rect 39858 136102 40478 136170
rect 39858 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 40478 136102
rect 39858 135978 40478 136046
rect 39858 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 40478 135978
rect 39858 118350 40478 135922
rect 61106 130350 61582 130384
rect 61106 130294 61130 130350
rect 61186 130294 61254 130350
rect 61310 130294 61378 130350
rect 61434 130294 61502 130350
rect 61558 130294 61582 130350
rect 61106 130226 61582 130294
rect 61106 130170 61130 130226
rect 61186 130170 61254 130226
rect 61310 130170 61378 130226
rect 61434 130170 61502 130226
rect 61558 130170 61582 130226
rect 61106 130102 61582 130170
rect 61106 130046 61130 130102
rect 61186 130046 61254 130102
rect 61310 130046 61378 130102
rect 61434 130046 61502 130102
rect 61558 130046 61582 130102
rect 61106 129978 61582 130046
rect 61106 129922 61130 129978
rect 61186 129922 61254 129978
rect 61310 129922 61378 129978
rect 61434 129922 61502 129978
rect 61558 129922 61582 129978
rect 61106 129888 61582 129922
rect 66858 130350 67478 147922
rect 66858 130294 66954 130350
rect 67010 130294 67078 130350
rect 67134 130294 67202 130350
rect 67258 130294 67326 130350
rect 67382 130294 67478 130350
rect 66858 130226 67478 130294
rect 66858 130170 66954 130226
rect 67010 130170 67078 130226
rect 67134 130170 67202 130226
rect 67258 130170 67326 130226
rect 67382 130170 67478 130226
rect 66858 130102 67478 130170
rect 66858 130046 66954 130102
rect 67010 130046 67078 130102
rect 67134 130046 67202 130102
rect 67258 130046 67326 130102
rect 67382 130046 67478 130102
rect 66858 129978 67478 130046
rect 66858 129922 66954 129978
rect 67010 129922 67078 129978
rect 67134 129922 67202 129978
rect 67258 129922 67326 129978
rect 67382 129922 67478 129978
rect 39858 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 40478 118350
rect 39858 118226 40478 118294
rect 39858 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 40478 118226
rect 39858 118102 40478 118170
rect 39858 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 40478 118102
rect 39858 117978 40478 118046
rect 39858 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 40478 117978
rect 39858 100350 40478 117922
rect 61906 118350 62382 118384
rect 61906 118294 61930 118350
rect 61986 118294 62054 118350
rect 62110 118294 62178 118350
rect 62234 118294 62302 118350
rect 62358 118294 62382 118350
rect 61906 118226 62382 118294
rect 61906 118170 61930 118226
rect 61986 118170 62054 118226
rect 62110 118170 62178 118226
rect 62234 118170 62302 118226
rect 62358 118170 62382 118226
rect 61906 118102 62382 118170
rect 61906 118046 61930 118102
rect 61986 118046 62054 118102
rect 62110 118046 62178 118102
rect 62234 118046 62302 118102
rect 62358 118046 62382 118102
rect 61906 117978 62382 118046
rect 61906 117922 61930 117978
rect 61986 117922 62054 117978
rect 62110 117922 62178 117978
rect 62234 117922 62302 117978
rect 62358 117922 62382 117978
rect 61906 117888 62382 117922
rect 61106 112350 61582 112384
rect 61106 112294 61130 112350
rect 61186 112294 61254 112350
rect 61310 112294 61378 112350
rect 61434 112294 61502 112350
rect 61558 112294 61582 112350
rect 61106 112226 61582 112294
rect 61106 112170 61130 112226
rect 61186 112170 61254 112226
rect 61310 112170 61378 112226
rect 61434 112170 61502 112226
rect 61558 112170 61582 112226
rect 61106 112102 61582 112170
rect 61106 112046 61130 112102
rect 61186 112046 61254 112102
rect 61310 112046 61378 112102
rect 61434 112046 61502 112102
rect 61558 112046 61582 112102
rect 61106 111978 61582 112046
rect 61106 111922 61130 111978
rect 61186 111922 61254 111978
rect 61310 111922 61378 111978
rect 61434 111922 61502 111978
rect 61558 111922 61582 111978
rect 61106 111888 61582 111922
rect 66858 112350 67478 129922
rect 66858 112294 66954 112350
rect 67010 112294 67078 112350
rect 67134 112294 67202 112350
rect 67258 112294 67326 112350
rect 67382 112294 67478 112350
rect 66858 112226 67478 112294
rect 66858 112170 66954 112226
rect 67010 112170 67078 112226
rect 67134 112170 67202 112226
rect 67258 112170 67326 112226
rect 67382 112170 67478 112226
rect 66858 112102 67478 112170
rect 66858 112046 66954 112102
rect 67010 112046 67078 112102
rect 67134 112046 67202 112102
rect 67258 112046 67326 112102
rect 67382 112046 67478 112102
rect 66858 111978 67478 112046
rect 66858 111922 66954 111978
rect 67010 111922 67078 111978
rect 67134 111922 67202 111978
rect 67258 111922 67326 111978
rect 67382 111922 67478 111978
rect 39858 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 40478 100350
rect 39858 100226 40478 100294
rect 39858 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 40478 100226
rect 39858 100102 40478 100170
rect 39858 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 40478 100102
rect 39858 99978 40478 100046
rect 39858 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 40478 99978
rect 39858 82350 40478 99922
rect 61906 100350 62382 100384
rect 61906 100294 61930 100350
rect 61986 100294 62054 100350
rect 62110 100294 62178 100350
rect 62234 100294 62302 100350
rect 62358 100294 62382 100350
rect 61906 100226 62382 100294
rect 61906 100170 61930 100226
rect 61986 100170 62054 100226
rect 62110 100170 62178 100226
rect 62234 100170 62302 100226
rect 62358 100170 62382 100226
rect 61906 100102 62382 100170
rect 61906 100046 61930 100102
rect 61986 100046 62054 100102
rect 62110 100046 62178 100102
rect 62234 100046 62302 100102
rect 62358 100046 62382 100102
rect 61906 99978 62382 100046
rect 61906 99922 61930 99978
rect 61986 99922 62054 99978
rect 62110 99922 62178 99978
rect 62234 99922 62302 99978
rect 62358 99922 62382 99978
rect 61906 99888 62382 99922
rect 61106 94350 61582 94384
rect 61106 94294 61130 94350
rect 61186 94294 61254 94350
rect 61310 94294 61378 94350
rect 61434 94294 61502 94350
rect 61558 94294 61582 94350
rect 61106 94226 61582 94294
rect 61106 94170 61130 94226
rect 61186 94170 61254 94226
rect 61310 94170 61378 94226
rect 61434 94170 61502 94226
rect 61558 94170 61582 94226
rect 61106 94102 61582 94170
rect 61106 94046 61130 94102
rect 61186 94046 61254 94102
rect 61310 94046 61378 94102
rect 61434 94046 61502 94102
rect 61558 94046 61582 94102
rect 61106 93978 61582 94046
rect 61106 93922 61130 93978
rect 61186 93922 61254 93978
rect 61310 93922 61378 93978
rect 61434 93922 61502 93978
rect 61558 93922 61582 93978
rect 61106 93888 61582 93922
rect 66858 94350 67478 111922
rect 66858 94294 66954 94350
rect 67010 94294 67078 94350
rect 67134 94294 67202 94350
rect 67258 94294 67326 94350
rect 67382 94294 67478 94350
rect 66858 94226 67478 94294
rect 66858 94170 66954 94226
rect 67010 94170 67078 94226
rect 67134 94170 67202 94226
rect 67258 94170 67326 94226
rect 67382 94170 67478 94226
rect 66858 94102 67478 94170
rect 66858 94046 66954 94102
rect 67010 94046 67078 94102
rect 67134 94046 67202 94102
rect 67258 94046 67326 94102
rect 67382 94046 67478 94102
rect 66858 93978 67478 94046
rect 66858 93922 66954 93978
rect 67010 93922 67078 93978
rect 67134 93922 67202 93978
rect 67258 93922 67326 93978
rect 67382 93922 67478 93978
rect 39858 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 40478 82350
rect 39858 82226 40478 82294
rect 39858 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 40478 82226
rect 39858 82102 40478 82170
rect 39858 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 40478 82102
rect 39858 81978 40478 82046
rect 39858 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 40478 81978
rect 39858 64350 40478 81922
rect 61906 82350 62382 82384
rect 61906 82294 61930 82350
rect 61986 82294 62054 82350
rect 62110 82294 62178 82350
rect 62234 82294 62302 82350
rect 62358 82294 62382 82350
rect 61906 82226 62382 82294
rect 61906 82170 61930 82226
rect 61986 82170 62054 82226
rect 62110 82170 62178 82226
rect 62234 82170 62302 82226
rect 62358 82170 62382 82226
rect 61906 82102 62382 82170
rect 61906 82046 61930 82102
rect 61986 82046 62054 82102
rect 62110 82046 62178 82102
rect 62234 82046 62302 82102
rect 62358 82046 62382 82102
rect 61906 81978 62382 82046
rect 61906 81922 61930 81978
rect 61986 81922 62054 81978
rect 62110 81922 62178 81978
rect 62234 81922 62302 81978
rect 62358 81922 62382 81978
rect 61906 81888 62382 81922
rect 61106 76350 61582 76384
rect 61106 76294 61130 76350
rect 61186 76294 61254 76350
rect 61310 76294 61378 76350
rect 61434 76294 61502 76350
rect 61558 76294 61582 76350
rect 61106 76226 61582 76294
rect 61106 76170 61130 76226
rect 61186 76170 61254 76226
rect 61310 76170 61378 76226
rect 61434 76170 61502 76226
rect 61558 76170 61582 76226
rect 61106 76102 61582 76170
rect 61106 76046 61130 76102
rect 61186 76046 61254 76102
rect 61310 76046 61378 76102
rect 61434 76046 61502 76102
rect 61558 76046 61582 76102
rect 61106 75978 61582 76046
rect 61106 75922 61130 75978
rect 61186 75922 61254 75978
rect 61310 75922 61378 75978
rect 61434 75922 61502 75978
rect 61558 75922 61582 75978
rect 61106 75888 61582 75922
rect 66858 76350 67478 93922
rect 66858 76294 66954 76350
rect 67010 76294 67078 76350
rect 67134 76294 67202 76350
rect 67258 76294 67326 76350
rect 67382 76294 67478 76350
rect 66858 76226 67478 76294
rect 66858 76170 66954 76226
rect 67010 76170 67078 76226
rect 67134 76170 67202 76226
rect 67258 76170 67326 76226
rect 67382 76170 67478 76226
rect 66858 76102 67478 76170
rect 66858 76046 66954 76102
rect 67010 76046 67078 76102
rect 67134 76046 67202 76102
rect 67258 76046 67326 76102
rect 67382 76046 67478 76102
rect 66858 75978 67478 76046
rect 66858 75922 66954 75978
rect 67010 75922 67078 75978
rect 67134 75922 67202 75978
rect 67258 75922 67326 75978
rect 67382 75922 67478 75978
rect 39858 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 40478 64350
rect 39858 64226 40478 64294
rect 39858 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 40478 64226
rect 39858 64102 40478 64170
rect 39858 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 40478 64102
rect 39858 63978 40478 64046
rect 39858 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 40478 63978
rect 39858 46350 40478 63922
rect 61906 64350 62382 64384
rect 61906 64294 61930 64350
rect 61986 64294 62054 64350
rect 62110 64294 62178 64350
rect 62234 64294 62302 64350
rect 62358 64294 62382 64350
rect 61906 64226 62382 64294
rect 61906 64170 61930 64226
rect 61986 64170 62054 64226
rect 62110 64170 62178 64226
rect 62234 64170 62302 64226
rect 62358 64170 62382 64226
rect 61906 64102 62382 64170
rect 61906 64046 61930 64102
rect 61986 64046 62054 64102
rect 62110 64046 62178 64102
rect 62234 64046 62302 64102
rect 62358 64046 62382 64102
rect 61906 63978 62382 64046
rect 61906 63922 61930 63978
rect 61986 63922 62054 63978
rect 62110 63922 62178 63978
rect 62234 63922 62302 63978
rect 62358 63922 62382 63978
rect 61906 63888 62382 63922
rect 61106 58350 61582 58384
rect 61106 58294 61130 58350
rect 61186 58294 61254 58350
rect 61310 58294 61378 58350
rect 61434 58294 61502 58350
rect 61558 58294 61582 58350
rect 61106 58226 61582 58294
rect 61106 58170 61130 58226
rect 61186 58170 61254 58226
rect 61310 58170 61378 58226
rect 61434 58170 61502 58226
rect 61558 58170 61582 58226
rect 61106 58102 61582 58170
rect 61106 58046 61130 58102
rect 61186 58046 61254 58102
rect 61310 58046 61378 58102
rect 61434 58046 61502 58102
rect 61558 58046 61582 58102
rect 61106 57978 61582 58046
rect 61106 57922 61130 57978
rect 61186 57922 61254 57978
rect 61310 57922 61378 57978
rect 61434 57922 61502 57978
rect 61558 57922 61582 57978
rect 61106 57888 61582 57922
rect 66858 58350 67478 75922
rect 66858 58294 66954 58350
rect 67010 58294 67078 58350
rect 67134 58294 67202 58350
rect 67258 58294 67326 58350
rect 67382 58294 67478 58350
rect 66858 58226 67478 58294
rect 66858 58170 66954 58226
rect 67010 58170 67078 58226
rect 67134 58170 67202 58226
rect 67258 58170 67326 58226
rect 67382 58170 67478 58226
rect 66858 58102 67478 58170
rect 66858 58046 66954 58102
rect 67010 58046 67078 58102
rect 67134 58046 67202 58102
rect 67258 58046 67326 58102
rect 67382 58046 67478 58102
rect 66858 57978 67478 58046
rect 66858 57922 66954 57978
rect 67010 57922 67078 57978
rect 67134 57922 67202 57978
rect 67258 57922 67326 57978
rect 67382 57922 67478 57978
rect 39858 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 40478 46350
rect 39858 46226 40478 46294
rect 39858 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 40478 46226
rect 39858 46102 40478 46170
rect 39858 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 40478 46102
rect 39858 45978 40478 46046
rect 39858 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 40478 45978
rect 39858 28350 40478 45922
rect 61906 46350 62382 46384
rect 61906 46294 61930 46350
rect 61986 46294 62054 46350
rect 62110 46294 62178 46350
rect 62234 46294 62302 46350
rect 62358 46294 62382 46350
rect 61906 46226 62382 46294
rect 61906 46170 61930 46226
rect 61986 46170 62054 46226
rect 62110 46170 62178 46226
rect 62234 46170 62302 46226
rect 62358 46170 62382 46226
rect 61906 46102 62382 46170
rect 61906 46046 61930 46102
rect 61986 46046 62054 46102
rect 62110 46046 62178 46102
rect 62234 46046 62302 46102
rect 62358 46046 62382 46102
rect 61906 45978 62382 46046
rect 61906 45922 61930 45978
rect 61986 45922 62054 45978
rect 62110 45922 62178 45978
rect 62234 45922 62302 45978
rect 62358 45922 62382 45978
rect 61906 45888 62382 45922
rect 39858 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 40478 28350
rect 39858 28226 40478 28294
rect 39858 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 40478 28226
rect 39858 28102 40478 28170
rect 39858 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 40478 28102
rect 39858 27978 40478 28046
rect 39858 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 40478 27978
rect 39858 10350 40478 27922
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 39858 -1120 40478 9922
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 40350 67478 57922
rect 66858 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 67478 40350
rect 66858 40226 67478 40294
rect 66858 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 67478 40226
rect 66858 40102 67478 40170
rect 66858 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 67478 40102
rect 66858 39978 67478 40046
rect 66858 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 67478 39978
rect 66858 22350 67478 39922
rect 66858 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 67478 22350
rect 66858 22226 67478 22294
rect 66858 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 67478 22226
rect 66858 22102 67478 22170
rect 66858 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 67478 22102
rect 66858 21978 67478 22046
rect 66858 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 67478 21978
rect 66858 4350 67478 21922
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 70364 227780 70420 227790
rect 70364 4228 70420 227724
rect 70364 4162 70420 4172
rect 70578 226350 71198 243922
rect 70578 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 71198 226350
rect 70578 226226 71198 226294
rect 70578 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 71198 226226
rect 70578 226102 71198 226170
rect 70578 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 71198 226102
rect 70578 225978 71198 226046
rect 70578 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 71198 225978
rect 70578 208350 71198 225922
rect 70578 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 71198 208350
rect 70578 208226 71198 208294
rect 70578 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 71198 208226
rect 70578 208102 71198 208170
rect 70578 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 71198 208102
rect 70578 207978 71198 208046
rect 70578 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 71198 207978
rect 70578 190350 71198 207922
rect 70578 190294 70674 190350
rect 70730 190294 70798 190350
rect 70854 190294 70922 190350
rect 70978 190294 71046 190350
rect 71102 190294 71198 190350
rect 70578 190226 71198 190294
rect 70578 190170 70674 190226
rect 70730 190170 70798 190226
rect 70854 190170 70922 190226
rect 70978 190170 71046 190226
rect 71102 190170 71198 190226
rect 70578 190102 71198 190170
rect 70578 190046 70674 190102
rect 70730 190046 70798 190102
rect 70854 190046 70922 190102
rect 70978 190046 71046 190102
rect 71102 190046 71198 190102
rect 70578 189978 71198 190046
rect 70578 189922 70674 189978
rect 70730 189922 70798 189978
rect 70854 189922 70922 189978
rect 70978 189922 71046 189978
rect 71102 189922 71198 189978
rect 70578 172350 71198 189922
rect 79808 190350 80128 190384
rect 79808 190294 79878 190350
rect 79934 190294 80002 190350
rect 80058 190294 80128 190350
rect 79808 190226 80128 190294
rect 79808 190170 79878 190226
rect 79934 190170 80002 190226
rect 80058 190170 80128 190226
rect 79808 190102 80128 190170
rect 79808 190046 79878 190102
rect 79934 190046 80002 190102
rect 80058 190046 80128 190102
rect 79808 189978 80128 190046
rect 79808 189922 79878 189978
rect 79934 189922 80002 189978
rect 80058 189922 80128 189978
rect 79808 189888 80128 189922
rect 70578 172294 70674 172350
rect 70730 172294 70798 172350
rect 70854 172294 70922 172350
rect 70978 172294 71046 172350
rect 71102 172294 71198 172350
rect 70578 172226 71198 172294
rect 70578 172170 70674 172226
rect 70730 172170 70798 172226
rect 70854 172170 70922 172226
rect 70978 172170 71046 172226
rect 71102 172170 71198 172226
rect 70578 172102 71198 172170
rect 70578 172046 70674 172102
rect 70730 172046 70798 172102
rect 70854 172046 70922 172102
rect 70978 172046 71046 172102
rect 71102 172046 71198 172102
rect 70578 171978 71198 172046
rect 70578 171922 70674 171978
rect 70730 171922 70798 171978
rect 70854 171922 70922 171978
rect 70978 171922 71046 171978
rect 71102 171922 71198 171978
rect 70578 154350 71198 171922
rect 79808 172350 80128 172384
rect 79808 172294 79878 172350
rect 79934 172294 80002 172350
rect 80058 172294 80128 172350
rect 79808 172226 80128 172294
rect 79808 172170 79878 172226
rect 79934 172170 80002 172226
rect 80058 172170 80128 172226
rect 79808 172102 80128 172170
rect 79808 172046 79878 172102
rect 79934 172046 80002 172102
rect 80058 172046 80128 172102
rect 79808 171978 80128 172046
rect 79808 171922 79878 171978
rect 79934 171922 80002 171978
rect 80058 171922 80128 171978
rect 79808 171888 80128 171922
rect 80556 158900 80612 158910
rect 70578 154294 70674 154350
rect 70730 154294 70798 154350
rect 70854 154294 70922 154350
rect 70978 154294 71046 154350
rect 71102 154294 71198 154350
rect 70578 154226 71198 154294
rect 70578 154170 70674 154226
rect 70730 154170 70798 154226
rect 70854 154170 70922 154226
rect 70978 154170 71046 154226
rect 71102 154170 71198 154226
rect 70578 154102 71198 154170
rect 70578 154046 70674 154102
rect 70730 154046 70798 154102
rect 70854 154046 70922 154102
rect 70978 154046 71046 154102
rect 71102 154046 71198 154102
rect 70578 153978 71198 154046
rect 70578 153922 70674 153978
rect 70730 153922 70798 153978
rect 70854 153922 70922 153978
rect 70978 153922 71046 153978
rect 71102 153922 71198 153978
rect 70578 136350 71198 153922
rect 70578 136294 70674 136350
rect 70730 136294 70798 136350
rect 70854 136294 70922 136350
rect 70978 136294 71046 136350
rect 71102 136294 71198 136350
rect 70578 136226 71198 136294
rect 70578 136170 70674 136226
rect 70730 136170 70798 136226
rect 70854 136170 70922 136226
rect 70978 136170 71046 136226
rect 71102 136170 71198 136226
rect 70578 136102 71198 136170
rect 70578 136046 70674 136102
rect 70730 136046 70798 136102
rect 70854 136046 70922 136102
rect 70978 136046 71046 136102
rect 71102 136046 71198 136102
rect 70578 135978 71198 136046
rect 70578 135922 70674 135978
rect 70730 135922 70798 135978
rect 70854 135922 70922 135978
rect 70978 135922 71046 135978
rect 71102 135922 71198 135978
rect 70578 118350 71198 135922
rect 70578 118294 70674 118350
rect 70730 118294 70798 118350
rect 70854 118294 70922 118350
rect 70978 118294 71046 118350
rect 71102 118294 71198 118350
rect 70578 118226 71198 118294
rect 70578 118170 70674 118226
rect 70730 118170 70798 118226
rect 70854 118170 70922 118226
rect 70978 118170 71046 118226
rect 71102 118170 71198 118226
rect 70578 118102 71198 118170
rect 70578 118046 70674 118102
rect 70730 118046 70798 118102
rect 70854 118046 70922 118102
rect 70978 118046 71046 118102
rect 71102 118046 71198 118102
rect 70578 117978 71198 118046
rect 70578 117922 70674 117978
rect 70730 117922 70798 117978
rect 70854 117922 70922 117978
rect 70978 117922 71046 117978
rect 71102 117922 71198 117978
rect 70578 100350 71198 117922
rect 70578 100294 70674 100350
rect 70730 100294 70798 100350
rect 70854 100294 70922 100350
rect 70978 100294 71046 100350
rect 71102 100294 71198 100350
rect 70578 100226 71198 100294
rect 70578 100170 70674 100226
rect 70730 100170 70798 100226
rect 70854 100170 70922 100226
rect 70978 100170 71046 100226
rect 71102 100170 71198 100226
rect 70578 100102 71198 100170
rect 70578 100046 70674 100102
rect 70730 100046 70798 100102
rect 70854 100046 70922 100102
rect 70978 100046 71046 100102
rect 71102 100046 71198 100102
rect 70578 99978 71198 100046
rect 70578 99922 70674 99978
rect 70730 99922 70798 99978
rect 70854 99922 70922 99978
rect 70978 99922 71046 99978
rect 71102 99922 71198 99978
rect 70578 82350 71198 99922
rect 70578 82294 70674 82350
rect 70730 82294 70798 82350
rect 70854 82294 70922 82350
rect 70978 82294 71046 82350
rect 71102 82294 71198 82350
rect 70578 82226 71198 82294
rect 70578 82170 70674 82226
rect 70730 82170 70798 82226
rect 70854 82170 70922 82226
rect 70978 82170 71046 82226
rect 71102 82170 71198 82226
rect 70578 82102 71198 82170
rect 70578 82046 70674 82102
rect 70730 82046 70798 82102
rect 70854 82046 70922 82102
rect 70978 82046 71046 82102
rect 71102 82046 71198 82102
rect 70578 81978 71198 82046
rect 70578 81922 70674 81978
rect 70730 81922 70798 81978
rect 70854 81922 70922 81978
rect 70978 81922 71046 81978
rect 71102 81922 71198 81978
rect 70578 64350 71198 81922
rect 70578 64294 70674 64350
rect 70730 64294 70798 64350
rect 70854 64294 70922 64350
rect 70978 64294 71046 64350
rect 71102 64294 71198 64350
rect 70578 64226 71198 64294
rect 70578 64170 70674 64226
rect 70730 64170 70798 64226
rect 70854 64170 70922 64226
rect 70978 64170 71046 64226
rect 71102 64170 71198 64226
rect 70578 64102 71198 64170
rect 70578 64046 70674 64102
rect 70730 64046 70798 64102
rect 70854 64046 70922 64102
rect 70978 64046 71046 64102
rect 71102 64046 71198 64102
rect 70578 63978 71198 64046
rect 70578 63922 70674 63978
rect 70730 63922 70798 63978
rect 70854 63922 70922 63978
rect 70978 63922 71046 63978
rect 71102 63922 71198 63978
rect 70578 46350 71198 63922
rect 70578 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 71198 46350
rect 70578 46226 71198 46294
rect 70578 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 71198 46226
rect 70578 46102 71198 46170
rect 70578 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 71198 46102
rect 70578 45978 71198 46046
rect 70578 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 71198 45978
rect 70578 28350 71198 45922
rect 70578 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 71198 28350
rect 70578 28226 71198 28294
rect 70578 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 71198 28226
rect 70578 28102 71198 28170
rect 70578 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 71198 28102
rect 70578 27978 71198 28046
rect 70578 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 71198 27978
rect 70578 10350 71198 27922
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 -1120 71198 9922
rect 78876 158788 78932 158798
rect 78876 4228 78932 158732
rect 78876 4162 78932 4172
rect 80556 4228 80612 158844
rect 81452 4340 81508 281372
rect 83132 280532 83188 374822
rect 83244 335998 83300 428428
rect 83580 427588 83636 427598
rect 83356 427476 83412 427486
rect 83356 408178 83412 427420
rect 83356 408112 83412 408122
rect 83468 425278 83524 425288
rect 83244 335932 83300 335942
rect 83356 374698 83412 374708
rect 83132 280466 83188 280476
rect 83356 280420 83412 374642
rect 83468 347698 83524 425222
rect 83580 409798 83636 427532
rect 97578 425262 98198 435922
rect 101298 478350 101918 493168
rect 101298 478294 101394 478350
rect 101450 478294 101518 478350
rect 101574 478294 101642 478350
rect 101698 478294 101766 478350
rect 101822 478294 101918 478350
rect 101298 478226 101918 478294
rect 101298 478170 101394 478226
rect 101450 478170 101518 478226
rect 101574 478170 101642 478226
rect 101698 478170 101766 478226
rect 101822 478170 101918 478226
rect 101298 478102 101918 478170
rect 101298 478046 101394 478102
rect 101450 478046 101518 478102
rect 101574 478046 101642 478102
rect 101698 478046 101766 478102
rect 101822 478046 101918 478102
rect 101298 477978 101918 478046
rect 101298 477922 101394 477978
rect 101450 477922 101518 477978
rect 101574 477922 101642 477978
rect 101698 477922 101766 477978
rect 101822 477922 101918 477978
rect 101298 460350 101918 477922
rect 101298 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 101918 460350
rect 101298 460226 101918 460294
rect 101298 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 101918 460226
rect 101298 460102 101918 460170
rect 101298 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 101918 460102
rect 101298 459978 101918 460046
rect 101298 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 101918 459978
rect 101298 442350 101918 459922
rect 101298 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 101918 442350
rect 101298 442226 101918 442294
rect 101298 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 101918 442226
rect 101298 442102 101918 442170
rect 101298 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 101918 442102
rect 101298 441978 101918 442046
rect 101298 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 101918 441978
rect 101298 425262 101918 441922
rect 121996 432628 122052 547982
rect 121996 432562 122052 432572
rect 128298 544350 128918 561922
rect 128298 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 128918 544350
rect 128298 544226 128918 544294
rect 128298 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 128918 544226
rect 128298 544102 128918 544170
rect 128298 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 128918 544102
rect 128298 543978 128918 544046
rect 128298 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 128918 543978
rect 128298 526350 128918 543922
rect 128298 526294 128394 526350
rect 128450 526294 128518 526350
rect 128574 526294 128642 526350
rect 128698 526294 128766 526350
rect 128822 526294 128918 526350
rect 128298 526226 128918 526294
rect 128298 526170 128394 526226
rect 128450 526170 128518 526226
rect 128574 526170 128642 526226
rect 128698 526170 128766 526226
rect 128822 526170 128918 526226
rect 128298 526102 128918 526170
rect 128298 526046 128394 526102
rect 128450 526046 128518 526102
rect 128574 526046 128642 526102
rect 128698 526046 128766 526102
rect 128822 526046 128918 526102
rect 128298 525978 128918 526046
rect 128298 525922 128394 525978
rect 128450 525922 128518 525978
rect 128574 525922 128642 525978
rect 128698 525922 128766 525978
rect 128822 525922 128918 525978
rect 128298 508350 128918 525922
rect 128298 508294 128394 508350
rect 128450 508294 128518 508350
rect 128574 508294 128642 508350
rect 128698 508294 128766 508350
rect 128822 508294 128918 508350
rect 128298 508226 128918 508294
rect 128298 508170 128394 508226
rect 128450 508170 128518 508226
rect 128574 508170 128642 508226
rect 128698 508170 128766 508226
rect 128822 508170 128918 508226
rect 128298 508102 128918 508170
rect 128298 508046 128394 508102
rect 128450 508046 128518 508102
rect 128574 508046 128642 508102
rect 128698 508046 128766 508102
rect 128822 508046 128918 508102
rect 128298 507978 128918 508046
rect 128298 507922 128394 507978
rect 128450 507922 128518 507978
rect 128574 507922 128642 507978
rect 128698 507922 128766 507978
rect 128822 507922 128918 507978
rect 128298 490350 128918 507922
rect 128298 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 128918 490350
rect 128298 490226 128918 490294
rect 128298 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 128918 490226
rect 128298 490102 128918 490170
rect 128298 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 128918 490102
rect 128298 489978 128918 490046
rect 128298 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 128918 489978
rect 128298 472350 128918 489922
rect 128298 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 128918 472350
rect 128298 472226 128918 472294
rect 128298 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 128918 472226
rect 128298 472102 128918 472170
rect 128298 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 128918 472102
rect 128298 471978 128918 472046
rect 128298 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 128918 471978
rect 128298 454350 128918 471922
rect 128298 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 128918 454350
rect 128298 454226 128918 454294
rect 128298 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 128918 454226
rect 128298 454102 128918 454170
rect 128298 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 128918 454102
rect 128298 453978 128918 454046
rect 128298 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 128918 453978
rect 128298 436350 128918 453922
rect 128298 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 128918 436350
rect 128298 436226 128918 436294
rect 128298 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 128918 436226
rect 128298 436102 128918 436170
rect 128298 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 128918 436102
rect 128298 435978 128918 436046
rect 128298 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 128918 435978
rect 128298 425262 128918 435922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 132018 568350 132638 585922
rect 132018 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 132638 568350
rect 132018 568226 132638 568294
rect 132018 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 132638 568226
rect 132018 568102 132638 568170
rect 132018 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 132638 568102
rect 132018 567978 132638 568046
rect 132018 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 132638 567978
rect 132018 550350 132638 567922
rect 132018 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 132638 550350
rect 132018 550226 132638 550294
rect 132018 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 132638 550226
rect 132018 550102 132638 550170
rect 132018 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 132638 550102
rect 132018 549978 132638 550046
rect 132018 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 132638 549978
rect 132018 532350 132638 549922
rect 132018 532294 132114 532350
rect 132170 532294 132238 532350
rect 132294 532294 132362 532350
rect 132418 532294 132486 532350
rect 132542 532294 132638 532350
rect 132018 532226 132638 532294
rect 132018 532170 132114 532226
rect 132170 532170 132238 532226
rect 132294 532170 132362 532226
rect 132418 532170 132486 532226
rect 132542 532170 132638 532226
rect 132018 532102 132638 532170
rect 132018 532046 132114 532102
rect 132170 532046 132238 532102
rect 132294 532046 132362 532102
rect 132418 532046 132486 532102
rect 132542 532046 132638 532102
rect 132018 531978 132638 532046
rect 132018 531922 132114 531978
rect 132170 531922 132238 531978
rect 132294 531922 132362 531978
rect 132418 531922 132486 531978
rect 132542 531922 132638 531978
rect 132018 514350 132638 531922
rect 132018 514294 132114 514350
rect 132170 514294 132238 514350
rect 132294 514294 132362 514350
rect 132418 514294 132486 514350
rect 132542 514294 132638 514350
rect 132018 514226 132638 514294
rect 132018 514170 132114 514226
rect 132170 514170 132238 514226
rect 132294 514170 132362 514226
rect 132418 514170 132486 514226
rect 132542 514170 132638 514226
rect 132018 514102 132638 514170
rect 132018 514046 132114 514102
rect 132170 514046 132238 514102
rect 132294 514046 132362 514102
rect 132418 514046 132486 514102
rect 132542 514046 132638 514102
rect 132018 513978 132638 514046
rect 132018 513922 132114 513978
rect 132170 513922 132238 513978
rect 132294 513922 132362 513978
rect 132418 513922 132486 513978
rect 132542 513922 132638 513978
rect 132018 496350 132638 513922
rect 132018 496294 132114 496350
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 132638 496350
rect 132018 496226 132638 496294
rect 132018 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 132638 496226
rect 132018 496102 132638 496170
rect 132018 496046 132114 496102
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 132638 496102
rect 132018 495978 132638 496046
rect 132018 495922 132114 495978
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 132638 495978
rect 132018 478350 132638 495922
rect 132018 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 132638 478350
rect 132018 478226 132638 478294
rect 132018 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 132638 478226
rect 132018 478102 132638 478170
rect 132018 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 132638 478102
rect 132018 477978 132638 478046
rect 132018 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 132638 477978
rect 132018 460350 132638 477922
rect 132018 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 132638 460350
rect 132018 460226 132638 460294
rect 132018 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 132638 460226
rect 132018 460102 132638 460170
rect 132018 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 132638 460102
rect 132018 459978 132638 460046
rect 132018 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 132638 459978
rect 132018 442350 132638 459922
rect 132018 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 132638 442350
rect 132018 442226 132638 442294
rect 132018 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 132638 442226
rect 132018 442102 132638 442170
rect 132018 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 132638 442102
rect 132018 441978 132638 442046
rect 132018 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 132638 441978
rect 132018 425262 132638 441922
rect 159018 597212 159638 598268
rect 159018 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 159638 597212
rect 159018 597088 159638 597156
rect 159018 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 159638 597088
rect 159018 596964 159638 597032
rect 159018 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 159638 596964
rect 159018 596840 159638 596908
rect 159018 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 159638 596840
rect 159018 580350 159638 596784
rect 159018 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 159638 580350
rect 159018 580226 159638 580294
rect 159018 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 159638 580226
rect 159018 580102 159638 580170
rect 159018 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 159638 580102
rect 159018 579978 159638 580046
rect 159018 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 159638 579978
rect 159018 562350 159638 579922
rect 159018 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 159638 562350
rect 159018 562226 159638 562294
rect 159018 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 159638 562226
rect 159018 562102 159638 562170
rect 159018 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 159638 562102
rect 159018 561978 159638 562046
rect 159018 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 159638 561978
rect 159018 544350 159638 561922
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 568350 163358 585922
rect 162738 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 163358 568350
rect 162738 568226 163358 568294
rect 162738 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 163358 568226
rect 162738 568102 163358 568170
rect 162738 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 163358 568102
rect 162738 567978 163358 568046
rect 162738 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 163358 567978
rect 162738 550350 163358 567922
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 189738 580350 190358 596784
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 189738 562350 190358 579922
rect 189738 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 190358 562350
rect 189738 562226 190358 562294
rect 189738 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 190358 562226
rect 189738 562102 190358 562170
rect 189738 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 190358 562102
rect 189738 561978 190358 562046
rect 189738 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 190358 561978
rect 162738 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 163358 550350
rect 162738 550226 163358 550294
rect 162738 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 163358 550226
rect 162738 550102 163358 550170
rect 162738 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 163358 550102
rect 162738 549978 163358 550046
rect 162738 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 163358 549978
rect 162738 548798 163358 549922
rect 179808 550350 180128 550384
rect 179808 550294 179878 550350
rect 179934 550294 180002 550350
rect 180058 550294 180128 550350
rect 179808 550226 180128 550294
rect 179808 550170 179878 550226
rect 179934 550170 180002 550226
rect 180058 550170 180128 550226
rect 179808 550102 180128 550170
rect 179808 550046 179878 550102
rect 179934 550046 180002 550102
rect 180058 550046 180128 550102
rect 179808 549978 180128 550046
rect 179808 549922 179878 549978
rect 179934 549922 180002 549978
rect 180058 549922 180128 549978
rect 179808 549888 180128 549922
rect 189738 548798 190358 561922
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 193458 586350 194078 597744
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 568350 194078 585922
rect 193458 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 194078 568350
rect 193458 568226 194078 568294
rect 193458 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 194078 568226
rect 193458 568102 194078 568170
rect 193458 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 194078 568102
rect 193458 567978 194078 568046
rect 193458 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 194078 567978
rect 193458 550350 194078 567922
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 220458 562350 221078 579922
rect 220458 562294 220554 562350
rect 220610 562294 220678 562350
rect 220734 562294 220802 562350
rect 220858 562294 220926 562350
rect 220982 562294 221078 562350
rect 220458 562226 221078 562294
rect 220458 562170 220554 562226
rect 220610 562170 220678 562226
rect 220734 562170 220802 562226
rect 220858 562170 220926 562226
rect 220982 562170 221078 562226
rect 220458 562102 221078 562170
rect 220458 562046 220554 562102
rect 220610 562046 220678 562102
rect 220734 562046 220802 562102
rect 220858 562046 220926 562102
rect 220982 562046 221078 562102
rect 220458 561978 221078 562046
rect 220458 561922 220554 561978
rect 220610 561922 220678 561978
rect 220734 561922 220802 561978
rect 220858 561922 220926 561978
rect 220982 561922 221078 561978
rect 212492 554372 212548 554382
rect 193458 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 194078 550350
rect 193458 550226 194078 550294
rect 193458 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 194078 550226
rect 193458 550102 194078 550170
rect 193458 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 194078 550102
rect 193458 549978 194078 550046
rect 193458 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 194078 549978
rect 193458 548798 194078 549922
rect 210528 550350 210848 550384
rect 210528 550294 210598 550350
rect 210654 550294 210722 550350
rect 210778 550294 210848 550350
rect 210528 550226 210848 550294
rect 210528 550170 210598 550226
rect 210654 550170 210722 550226
rect 210778 550170 210848 550226
rect 210528 550102 210848 550170
rect 210528 550046 210598 550102
rect 210654 550046 210722 550102
rect 210778 550046 210848 550102
rect 210528 549978 210848 550046
rect 210528 549922 210598 549978
rect 210654 549922 210722 549978
rect 210778 549922 210848 549978
rect 210528 549888 210848 549922
rect 159018 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 159638 544350
rect 159018 544226 159638 544294
rect 159018 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 159638 544226
rect 159018 544102 159638 544170
rect 159018 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 159638 544102
rect 159018 543978 159638 544046
rect 159018 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 159638 543978
rect 159018 526350 159638 543922
rect 164448 544350 164768 544384
rect 164448 544294 164518 544350
rect 164574 544294 164642 544350
rect 164698 544294 164768 544350
rect 164448 544226 164768 544294
rect 164448 544170 164518 544226
rect 164574 544170 164642 544226
rect 164698 544170 164768 544226
rect 164448 544102 164768 544170
rect 164448 544046 164518 544102
rect 164574 544046 164642 544102
rect 164698 544046 164768 544102
rect 164448 543978 164768 544046
rect 164448 543922 164518 543978
rect 164574 543922 164642 543978
rect 164698 543922 164768 543978
rect 164448 543888 164768 543922
rect 195168 544350 195488 544384
rect 195168 544294 195238 544350
rect 195294 544294 195362 544350
rect 195418 544294 195488 544350
rect 195168 544226 195488 544294
rect 195168 544170 195238 544226
rect 195294 544170 195362 544226
rect 195418 544170 195488 544226
rect 195168 544102 195488 544170
rect 195168 544046 195238 544102
rect 195294 544046 195362 544102
rect 195418 544046 195488 544102
rect 195168 543978 195488 544046
rect 195168 543922 195238 543978
rect 195294 543922 195362 543978
rect 195418 543922 195488 543978
rect 195168 543888 195488 543922
rect 179808 532350 180128 532384
rect 179808 532294 179878 532350
rect 179934 532294 180002 532350
rect 180058 532294 180128 532350
rect 179808 532226 180128 532294
rect 179808 532170 179878 532226
rect 179934 532170 180002 532226
rect 180058 532170 180128 532226
rect 179808 532102 180128 532170
rect 179808 532046 179878 532102
rect 179934 532046 180002 532102
rect 180058 532046 180128 532102
rect 179808 531978 180128 532046
rect 179808 531922 179878 531978
rect 179934 531922 180002 531978
rect 180058 531922 180128 531978
rect 179808 531888 180128 531922
rect 210528 532350 210848 532384
rect 210528 532294 210598 532350
rect 210654 532294 210722 532350
rect 210778 532294 210848 532350
rect 210528 532226 210848 532294
rect 210528 532170 210598 532226
rect 210654 532170 210722 532226
rect 210778 532170 210848 532226
rect 210528 532102 210848 532170
rect 210528 532046 210598 532102
rect 210654 532046 210722 532102
rect 210778 532046 210848 532102
rect 210528 531978 210848 532046
rect 210528 531922 210598 531978
rect 210654 531922 210722 531978
rect 210778 531922 210848 531978
rect 210528 531888 210848 531922
rect 159018 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 159638 526350
rect 159018 526226 159638 526294
rect 159018 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 159638 526226
rect 159018 526102 159638 526170
rect 159018 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 159638 526102
rect 159018 525978 159638 526046
rect 159018 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 159638 525978
rect 159018 508350 159638 525922
rect 164448 526350 164768 526384
rect 164448 526294 164518 526350
rect 164574 526294 164642 526350
rect 164698 526294 164768 526350
rect 164448 526226 164768 526294
rect 164448 526170 164518 526226
rect 164574 526170 164642 526226
rect 164698 526170 164768 526226
rect 164448 526102 164768 526170
rect 164448 526046 164518 526102
rect 164574 526046 164642 526102
rect 164698 526046 164768 526102
rect 164448 525978 164768 526046
rect 164448 525922 164518 525978
rect 164574 525922 164642 525978
rect 164698 525922 164768 525978
rect 164448 525888 164768 525922
rect 195168 526350 195488 526384
rect 195168 526294 195238 526350
rect 195294 526294 195362 526350
rect 195418 526294 195488 526350
rect 195168 526226 195488 526294
rect 195168 526170 195238 526226
rect 195294 526170 195362 526226
rect 195418 526170 195488 526226
rect 195168 526102 195488 526170
rect 195168 526046 195238 526102
rect 195294 526046 195362 526102
rect 195418 526046 195488 526102
rect 195168 525978 195488 526046
rect 195168 525922 195238 525978
rect 195294 525922 195362 525978
rect 195418 525922 195488 525978
rect 195168 525888 195488 525922
rect 179808 514350 180128 514384
rect 179808 514294 179878 514350
rect 179934 514294 180002 514350
rect 180058 514294 180128 514350
rect 179808 514226 180128 514294
rect 179808 514170 179878 514226
rect 179934 514170 180002 514226
rect 180058 514170 180128 514226
rect 179808 514102 180128 514170
rect 179808 514046 179878 514102
rect 179934 514046 180002 514102
rect 180058 514046 180128 514102
rect 179808 513978 180128 514046
rect 179808 513922 179878 513978
rect 179934 513922 180002 513978
rect 180058 513922 180128 513978
rect 179808 513888 180128 513922
rect 210528 514350 210848 514384
rect 210528 514294 210598 514350
rect 210654 514294 210722 514350
rect 210778 514294 210848 514350
rect 210528 514226 210848 514294
rect 210528 514170 210598 514226
rect 210654 514170 210722 514226
rect 210778 514170 210848 514226
rect 210528 514102 210848 514170
rect 210528 514046 210598 514102
rect 210654 514046 210722 514102
rect 210778 514046 210848 514102
rect 210528 513978 210848 514046
rect 210528 513922 210598 513978
rect 210654 513922 210722 513978
rect 210778 513922 210848 513978
rect 210528 513888 210848 513922
rect 159018 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 159638 508350
rect 159018 508226 159638 508294
rect 159018 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 159638 508226
rect 159018 508102 159638 508170
rect 159018 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 159638 508102
rect 159018 507978 159638 508046
rect 159018 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 159638 507978
rect 159018 490350 159638 507922
rect 164448 508350 164768 508384
rect 164448 508294 164518 508350
rect 164574 508294 164642 508350
rect 164698 508294 164768 508350
rect 164448 508226 164768 508294
rect 164448 508170 164518 508226
rect 164574 508170 164642 508226
rect 164698 508170 164768 508226
rect 164448 508102 164768 508170
rect 164448 508046 164518 508102
rect 164574 508046 164642 508102
rect 164698 508046 164768 508102
rect 164448 507978 164768 508046
rect 164448 507922 164518 507978
rect 164574 507922 164642 507978
rect 164698 507922 164768 507978
rect 164448 507888 164768 507922
rect 195168 508350 195488 508384
rect 195168 508294 195238 508350
rect 195294 508294 195362 508350
rect 195418 508294 195488 508350
rect 195168 508226 195488 508294
rect 195168 508170 195238 508226
rect 195294 508170 195362 508226
rect 195418 508170 195488 508226
rect 195168 508102 195488 508170
rect 195168 508046 195238 508102
rect 195294 508046 195362 508102
rect 195418 508046 195488 508102
rect 195168 507978 195488 508046
rect 195168 507922 195238 507978
rect 195294 507922 195362 507978
rect 195418 507922 195488 507978
rect 195168 507888 195488 507922
rect 176988 501732 177044 501742
rect 171500 501620 171556 501630
rect 159018 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 159638 490350
rect 159018 490226 159638 490294
rect 159018 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 159638 490226
rect 159018 490102 159638 490170
rect 159018 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 159638 490102
rect 159018 489978 159638 490046
rect 159018 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 159638 489978
rect 159018 472350 159638 489922
rect 159018 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 159638 472350
rect 159018 472226 159638 472294
rect 159018 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 159638 472226
rect 159018 472102 159638 472170
rect 159018 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 159638 472102
rect 159018 471978 159638 472046
rect 159018 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 159638 471978
rect 159018 454350 159638 471922
rect 159018 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 159638 454350
rect 159018 454226 159638 454294
rect 159018 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 159638 454226
rect 159018 454102 159638 454170
rect 159018 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 159638 454102
rect 159018 453978 159638 454046
rect 159018 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 159638 453978
rect 159018 436350 159638 453922
rect 159018 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 159638 436350
rect 159018 436226 159638 436294
rect 159018 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 159638 436226
rect 159018 436102 159638 436170
rect 159018 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 159638 436102
rect 159018 435978 159638 436046
rect 159018 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 159638 435978
rect 159018 425262 159638 435922
rect 162738 496350 163358 501266
rect 171500 500052 171556 501564
rect 176988 500612 177044 501676
rect 176988 500546 177044 500556
rect 171500 499986 171556 499996
rect 162738 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 163358 496350
rect 162738 496226 163358 496294
rect 162738 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 163358 496226
rect 162738 496102 163358 496170
rect 162738 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 163358 496102
rect 162738 495978 163358 496046
rect 162738 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 163358 495978
rect 162738 478350 163358 495922
rect 189738 490350 190358 501266
rect 189738 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 190358 490350
rect 189738 490226 190358 490294
rect 189738 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 190358 490226
rect 189738 490102 190358 490170
rect 189738 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 190358 490102
rect 189738 489978 190358 490046
rect 189738 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 190358 489978
rect 169596 488098 169652 488108
rect 162738 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 163358 478350
rect 162738 478226 163358 478294
rect 162738 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 163358 478226
rect 162738 478102 163358 478170
rect 162738 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 163358 478102
rect 162738 477978 163358 478046
rect 162738 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 163358 477978
rect 162738 460350 163358 477922
rect 166236 479638 166292 479648
rect 162738 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 163358 460350
rect 162738 460226 163358 460294
rect 162738 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 163358 460226
rect 162738 460102 163358 460170
rect 162738 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 163358 460102
rect 162738 459978 163358 460046
rect 162738 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 163358 459978
rect 162738 442350 163358 459922
rect 162738 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 163358 442350
rect 162738 442226 163358 442294
rect 162738 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 163358 442226
rect 162738 442102 163358 442170
rect 162738 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 163358 442102
rect 162738 441978 163358 442046
rect 162738 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 163358 441978
rect 162738 425262 163358 441922
rect 164556 472618 164612 472628
rect 164556 433412 164612 472562
rect 164556 433346 164612 433356
rect 166236 433412 166292 479582
rect 166236 433346 166292 433356
rect 169596 433412 169652 488042
rect 169596 433346 169652 433356
rect 189738 472350 190358 489922
rect 189738 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 190358 472350
rect 189738 472226 190358 472294
rect 189738 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 190358 472226
rect 189738 472102 190358 472170
rect 189738 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 190358 472102
rect 189738 471978 190358 472046
rect 189738 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 190358 471978
rect 189738 454350 190358 471922
rect 189738 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 190358 454350
rect 189738 454226 190358 454294
rect 189738 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 190358 454226
rect 189738 454102 190358 454170
rect 189738 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 190358 454102
rect 189738 453978 190358 454046
rect 189738 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 190358 453978
rect 189738 436350 190358 453922
rect 189738 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 190358 436350
rect 189738 436226 190358 436294
rect 189738 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 190358 436226
rect 189738 436102 190358 436170
rect 189738 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 190358 436102
rect 189738 435978 190358 436046
rect 189738 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 190358 435978
rect 189738 425262 190358 435922
rect 193458 496350 194078 501266
rect 193458 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 194078 496350
rect 193458 496226 194078 496294
rect 193458 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 194078 496226
rect 193458 496102 194078 496170
rect 193458 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 194078 496102
rect 193458 495978 194078 496046
rect 193458 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 194078 495978
rect 193458 478350 194078 495922
rect 193458 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 194078 478350
rect 193458 478226 194078 478294
rect 193458 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 194078 478226
rect 193458 478102 194078 478170
rect 193458 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 194078 478102
rect 193458 477978 194078 478046
rect 193458 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 194078 477978
rect 193458 460350 194078 477922
rect 193458 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 194078 460350
rect 193458 460226 194078 460294
rect 193458 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 194078 460226
rect 193458 460102 194078 460170
rect 193458 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 194078 460102
rect 193458 459978 194078 460046
rect 193458 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 194078 459978
rect 193458 442350 194078 459922
rect 193458 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 194078 442350
rect 193458 442226 194078 442294
rect 193458 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 194078 442226
rect 193458 442102 194078 442170
rect 193458 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 194078 442102
rect 193458 441978 194078 442046
rect 193458 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 194078 441978
rect 193458 425262 194078 441922
rect 212492 432740 212548 554316
rect 212492 430052 212548 432684
rect 212492 429986 212548 429996
rect 220458 544350 221078 561922
rect 220458 544294 220554 544350
rect 220610 544294 220678 544350
rect 220734 544294 220802 544350
rect 220858 544294 220926 544350
rect 220982 544294 221078 544350
rect 220458 544226 221078 544294
rect 220458 544170 220554 544226
rect 220610 544170 220678 544226
rect 220734 544170 220802 544226
rect 220858 544170 220926 544226
rect 220982 544170 221078 544226
rect 220458 544102 221078 544170
rect 220458 544046 220554 544102
rect 220610 544046 220678 544102
rect 220734 544046 220802 544102
rect 220858 544046 220926 544102
rect 220982 544046 221078 544102
rect 220458 543978 221078 544046
rect 220458 543922 220554 543978
rect 220610 543922 220678 543978
rect 220734 543922 220802 543978
rect 220858 543922 220926 543978
rect 220982 543922 221078 543978
rect 220458 526350 221078 543922
rect 220458 526294 220554 526350
rect 220610 526294 220678 526350
rect 220734 526294 220802 526350
rect 220858 526294 220926 526350
rect 220982 526294 221078 526350
rect 220458 526226 221078 526294
rect 220458 526170 220554 526226
rect 220610 526170 220678 526226
rect 220734 526170 220802 526226
rect 220858 526170 220926 526226
rect 220982 526170 221078 526226
rect 220458 526102 221078 526170
rect 220458 526046 220554 526102
rect 220610 526046 220678 526102
rect 220734 526046 220802 526102
rect 220858 526046 220926 526102
rect 220982 526046 221078 526102
rect 220458 525978 221078 526046
rect 220458 525922 220554 525978
rect 220610 525922 220678 525978
rect 220734 525922 220802 525978
rect 220858 525922 220926 525978
rect 220982 525922 221078 525978
rect 220458 508350 221078 525922
rect 220458 508294 220554 508350
rect 220610 508294 220678 508350
rect 220734 508294 220802 508350
rect 220858 508294 220926 508350
rect 220982 508294 221078 508350
rect 220458 508226 221078 508294
rect 220458 508170 220554 508226
rect 220610 508170 220678 508226
rect 220734 508170 220802 508226
rect 220858 508170 220926 508226
rect 220982 508170 221078 508226
rect 220458 508102 221078 508170
rect 220458 508046 220554 508102
rect 220610 508046 220678 508102
rect 220734 508046 220802 508102
rect 220858 508046 220926 508102
rect 220982 508046 221078 508102
rect 220458 507978 221078 508046
rect 220458 507922 220554 507978
rect 220610 507922 220678 507978
rect 220734 507922 220802 507978
rect 220858 507922 220926 507978
rect 220982 507922 221078 507978
rect 220458 490350 221078 507922
rect 220458 490294 220554 490350
rect 220610 490294 220678 490350
rect 220734 490294 220802 490350
rect 220858 490294 220926 490350
rect 220982 490294 221078 490350
rect 220458 490226 221078 490294
rect 220458 490170 220554 490226
rect 220610 490170 220678 490226
rect 220734 490170 220802 490226
rect 220858 490170 220926 490226
rect 220982 490170 221078 490226
rect 220458 490102 221078 490170
rect 220458 490046 220554 490102
rect 220610 490046 220678 490102
rect 220734 490046 220802 490102
rect 220858 490046 220926 490102
rect 220982 490046 221078 490102
rect 220458 489978 221078 490046
rect 220458 489922 220554 489978
rect 220610 489922 220678 489978
rect 220734 489922 220802 489978
rect 220858 489922 220926 489978
rect 220982 489922 221078 489978
rect 220458 472350 221078 489922
rect 220458 472294 220554 472350
rect 220610 472294 220678 472350
rect 220734 472294 220802 472350
rect 220858 472294 220926 472350
rect 220982 472294 221078 472350
rect 220458 472226 221078 472294
rect 220458 472170 220554 472226
rect 220610 472170 220678 472226
rect 220734 472170 220802 472226
rect 220858 472170 220926 472226
rect 220982 472170 221078 472226
rect 220458 472102 221078 472170
rect 220458 472046 220554 472102
rect 220610 472046 220678 472102
rect 220734 472046 220802 472102
rect 220858 472046 220926 472102
rect 220982 472046 221078 472102
rect 220458 471978 221078 472046
rect 220458 471922 220554 471978
rect 220610 471922 220678 471978
rect 220734 471922 220802 471978
rect 220858 471922 220926 471978
rect 220982 471922 221078 471978
rect 220458 454350 221078 471922
rect 220458 454294 220554 454350
rect 220610 454294 220678 454350
rect 220734 454294 220802 454350
rect 220858 454294 220926 454350
rect 220982 454294 221078 454350
rect 220458 454226 221078 454294
rect 220458 454170 220554 454226
rect 220610 454170 220678 454226
rect 220734 454170 220802 454226
rect 220858 454170 220926 454226
rect 220982 454170 221078 454226
rect 220458 454102 221078 454170
rect 220458 454046 220554 454102
rect 220610 454046 220678 454102
rect 220734 454046 220802 454102
rect 220858 454046 220926 454102
rect 220982 454046 221078 454102
rect 220458 453978 221078 454046
rect 220458 453922 220554 453978
rect 220610 453922 220678 453978
rect 220734 453922 220802 453978
rect 220858 453922 220926 453978
rect 220982 453922 221078 453978
rect 220458 436350 221078 453922
rect 220458 436294 220554 436350
rect 220610 436294 220678 436350
rect 220734 436294 220802 436350
rect 220858 436294 220926 436350
rect 220982 436294 221078 436350
rect 220458 436226 221078 436294
rect 220458 436170 220554 436226
rect 220610 436170 220678 436226
rect 220734 436170 220802 436226
rect 220858 436170 220926 436226
rect 220982 436170 221078 436226
rect 220458 436102 221078 436170
rect 220458 436046 220554 436102
rect 220610 436046 220678 436102
rect 220734 436046 220802 436102
rect 220858 436046 220926 436102
rect 220982 436046 221078 436102
rect 220458 435978 221078 436046
rect 220458 435922 220554 435978
rect 220610 435922 220678 435978
rect 220734 435922 220802 435978
rect 220858 435922 220926 435978
rect 220982 435922 221078 435978
rect 220458 425262 221078 435922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 568350 224798 585922
rect 224178 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 224798 568350
rect 224178 568226 224798 568294
rect 224178 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 224798 568226
rect 224178 568102 224798 568170
rect 224178 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 224798 568102
rect 224178 567978 224798 568046
rect 224178 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 224798 567978
rect 224178 550350 224798 567922
rect 224178 550294 224274 550350
rect 224330 550294 224398 550350
rect 224454 550294 224522 550350
rect 224578 550294 224646 550350
rect 224702 550294 224798 550350
rect 224178 550226 224798 550294
rect 224178 550170 224274 550226
rect 224330 550170 224398 550226
rect 224454 550170 224522 550226
rect 224578 550170 224646 550226
rect 224702 550170 224798 550226
rect 224178 550102 224798 550170
rect 224178 550046 224274 550102
rect 224330 550046 224398 550102
rect 224454 550046 224522 550102
rect 224578 550046 224646 550102
rect 224702 550046 224798 550102
rect 224178 549978 224798 550046
rect 224178 549922 224274 549978
rect 224330 549922 224398 549978
rect 224454 549922 224522 549978
rect 224578 549922 224646 549978
rect 224702 549922 224798 549978
rect 224178 532350 224798 549922
rect 224178 532294 224274 532350
rect 224330 532294 224398 532350
rect 224454 532294 224522 532350
rect 224578 532294 224646 532350
rect 224702 532294 224798 532350
rect 224178 532226 224798 532294
rect 224178 532170 224274 532226
rect 224330 532170 224398 532226
rect 224454 532170 224522 532226
rect 224578 532170 224646 532226
rect 224702 532170 224798 532226
rect 224178 532102 224798 532170
rect 224178 532046 224274 532102
rect 224330 532046 224398 532102
rect 224454 532046 224522 532102
rect 224578 532046 224646 532102
rect 224702 532046 224798 532102
rect 224178 531978 224798 532046
rect 224178 531922 224274 531978
rect 224330 531922 224398 531978
rect 224454 531922 224522 531978
rect 224578 531922 224646 531978
rect 224702 531922 224798 531978
rect 224178 514350 224798 531922
rect 224178 514294 224274 514350
rect 224330 514294 224398 514350
rect 224454 514294 224522 514350
rect 224578 514294 224646 514350
rect 224702 514294 224798 514350
rect 224178 514226 224798 514294
rect 224178 514170 224274 514226
rect 224330 514170 224398 514226
rect 224454 514170 224522 514226
rect 224578 514170 224646 514226
rect 224702 514170 224798 514226
rect 224178 514102 224798 514170
rect 224178 514046 224274 514102
rect 224330 514046 224398 514102
rect 224454 514046 224522 514102
rect 224578 514046 224646 514102
rect 224702 514046 224798 514102
rect 224178 513978 224798 514046
rect 224178 513922 224274 513978
rect 224330 513922 224398 513978
rect 224454 513922 224522 513978
rect 224578 513922 224646 513978
rect 224702 513922 224798 513978
rect 224178 496350 224798 513922
rect 224178 496294 224274 496350
rect 224330 496294 224398 496350
rect 224454 496294 224522 496350
rect 224578 496294 224646 496350
rect 224702 496294 224798 496350
rect 224178 496226 224798 496294
rect 224178 496170 224274 496226
rect 224330 496170 224398 496226
rect 224454 496170 224522 496226
rect 224578 496170 224646 496226
rect 224702 496170 224798 496226
rect 224178 496102 224798 496170
rect 224178 496046 224274 496102
rect 224330 496046 224398 496102
rect 224454 496046 224522 496102
rect 224578 496046 224646 496102
rect 224702 496046 224798 496102
rect 224178 495978 224798 496046
rect 224178 495922 224274 495978
rect 224330 495922 224398 495978
rect 224454 495922 224522 495978
rect 224578 495922 224646 495978
rect 224702 495922 224798 495978
rect 224178 478350 224798 495922
rect 224178 478294 224274 478350
rect 224330 478294 224398 478350
rect 224454 478294 224522 478350
rect 224578 478294 224646 478350
rect 224702 478294 224798 478350
rect 224178 478226 224798 478294
rect 224178 478170 224274 478226
rect 224330 478170 224398 478226
rect 224454 478170 224522 478226
rect 224578 478170 224646 478226
rect 224702 478170 224798 478226
rect 224178 478102 224798 478170
rect 224178 478046 224274 478102
rect 224330 478046 224398 478102
rect 224454 478046 224522 478102
rect 224578 478046 224646 478102
rect 224702 478046 224798 478102
rect 224178 477978 224798 478046
rect 224178 477922 224274 477978
rect 224330 477922 224398 477978
rect 224454 477922 224522 477978
rect 224578 477922 224646 477978
rect 224702 477922 224798 477978
rect 224178 460350 224798 477922
rect 224178 460294 224274 460350
rect 224330 460294 224398 460350
rect 224454 460294 224522 460350
rect 224578 460294 224646 460350
rect 224702 460294 224798 460350
rect 224178 460226 224798 460294
rect 224178 460170 224274 460226
rect 224330 460170 224398 460226
rect 224454 460170 224522 460226
rect 224578 460170 224646 460226
rect 224702 460170 224798 460226
rect 224178 460102 224798 460170
rect 224178 460046 224274 460102
rect 224330 460046 224398 460102
rect 224454 460046 224522 460102
rect 224578 460046 224646 460102
rect 224702 460046 224798 460102
rect 224178 459978 224798 460046
rect 224178 459922 224274 459978
rect 224330 459922 224398 459978
rect 224454 459922 224522 459978
rect 224578 459922 224646 459978
rect 224702 459922 224798 459978
rect 224178 442350 224798 459922
rect 224178 442294 224274 442350
rect 224330 442294 224398 442350
rect 224454 442294 224522 442350
rect 224578 442294 224646 442350
rect 224702 442294 224798 442350
rect 224178 442226 224798 442294
rect 224178 442170 224274 442226
rect 224330 442170 224398 442226
rect 224454 442170 224522 442226
rect 224578 442170 224646 442226
rect 224702 442170 224798 442226
rect 224178 442102 224798 442170
rect 224178 442046 224274 442102
rect 224330 442046 224398 442102
rect 224454 442046 224522 442102
rect 224578 442046 224646 442102
rect 224702 442046 224798 442102
rect 224178 441978 224798 442046
rect 224178 441922 224274 441978
rect 224330 441922 224398 441978
rect 224454 441922 224522 441978
rect 224578 441922 224646 441978
rect 224702 441922 224798 441978
rect 224178 425262 224798 441922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 251178 562350 251798 579922
rect 251178 562294 251274 562350
rect 251330 562294 251398 562350
rect 251454 562294 251522 562350
rect 251578 562294 251646 562350
rect 251702 562294 251798 562350
rect 251178 562226 251798 562294
rect 251178 562170 251274 562226
rect 251330 562170 251398 562226
rect 251454 562170 251522 562226
rect 251578 562170 251646 562226
rect 251702 562170 251798 562226
rect 251178 562102 251798 562170
rect 251178 562046 251274 562102
rect 251330 562046 251398 562102
rect 251454 562046 251522 562102
rect 251578 562046 251646 562102
rect 251702 562046 251798 562102
rect 251178 561978 251798 562046
rect 251178 561922 251274 561978
rect 251330 561922 251398 561978
rect 251454 561922 251522 561978
rect 251578 561922 251646 561978
rect 251702 561922 251798 561978
rect 251178 544350 251798 561922
rect 251178 544294 251274 544350
rect 251330 544294 251398 544350
rect 251454 544294 251522 544350
rect 251578 544294 251646 544350
rect 251702 544294 251798 544350
rect 251178 544226 251798 544294
rect 251178 544170 251274 544226
rect 251330 544170 251398 544226
rect 251454 544170 251522 544226
rect 251578 544170 251646 544226
rect 251702 544170 251798 544226
rect 251178 544102 251798 544170
rect 251178 544046 251274 544102
rect 251330 544046 251398 544102
rect 251454 544046 251522 544102
rect 251578 544046 251646 544102
rect 251702 544046 251798 544102
rect 251178 543978 251798 544046
rect 251178 543922 251274 543978
rect 251330 543922 251398 543978
rect 251454 543922 251522 543978
rect 251578 543922 251646 543978
rect 251702 543922 251798 543978
rect 251178 526350 251798 543922
rect 251178 526294 251274 526350
rect 251330 526294 251398 526350
rect 251454 526294 251522 526350
rect 251578 526294 251646 526350
rect 251702 526294 251798 526350
rect 251178 526226 251798 526294
rect 251178 526170 251274 526226
rect 251330 526170 251398 526226
rect 251454 526170 251522 526226
rect 251578 526170 251646 526226
rect 251702 526170 251798 526226
rect 251178 526102 251798 526170
rect 251178 526046 251274 526102
rect 251330 526046 251398 526102
rect 251454 526046 251522 526102
rect 251578 526046 251646 526102
rect 251702 526046 251798 526102
rect 251178 525978 251798 526046
rect 251178 525922 251274 525978
rect 251330 525922 251398 525978
rect 251454 525922 251522 525978
rect 251578 525922 251646 525978
rect 251702 525922 251798 525978
rect 251178 508350 251798 525922
rect 251178 508294 251274 508350
rect 251330 508294 251398 508350
rect 251454 508294 251522 508350
rect 251578 508294 251646 508350
rect 251702 508294 251798 508350
rect 251178 508226 251798 508294
rect 251178 508170 251274 508226
rect 251330 508170 251398 508226
rect 251454 508170 251522 508226
rect 251578 508170 251646 508226
rect 251702 508170 251798 508226
rect 251178 508102 251798 508170
rect 251178 508046 251274 508102
rect 251330 508046 251398 508102
rect 251454 508046 251522 508102
rect 251578 508046 251646 508102
rect 251702 508046 251798 508102
rect 251178 507978 251798 508046
rect 251178 507922 251274 507978
rect 251330 507922 251398 507978
rect 251454 507922 251522 507978
rect 251578 507922 251646 507978
rect 251702 507922 251798 507978
rect 251178 490350 251798 507922
rect 251178 490294 251274 490350
rect 251330 490294 251398 490350
rect 251454 490294 251522 490350
rect 251578 490294 251646 490350
rect 251702 490294 251798 490350
rect 251178 490226 251798 490294
rect 251178 490170 251274 490226
rect 251330 490170 251398 490226
rect 251454 490170 251522 490226
rect 251578 490170 251646 490226
rect 251702 490170 251798 490226
rect 251178 490102 251798 490170
rect 251178 490046 251274 490102
rect 251330 490046 251398 490102
rect 251454 490046 251522 490102
rect 251578 490046 251646 490102
rect 251702 490046 251798 490102
rect 251178 489978 251798 490046
rect 251178 489922 251274 489978
rect 251330 489922 251398 489978
rect 251454 489922 251522 489978
rect 251578 489922 251646 489978
rect 251702 489922 251798 489978
rect 251178 472350 251798 489922
rect 251178 472294 251274 472350
rect 251330 472294 251398 472350
rect 251454 472294 251522 472350
rect 251578 472294 251646 472350
rect 251702 472294 251798 472350
rect 251178 472226 251798 472294
rect 251178 472170 251274 472226
rect 251330 472170 251398 472226
rect 251454 472170 251522 472226
rect 251578 472170 251646 472226
rect 251702 472170 251798 472226
rect 251178 472102 251798 472170
rect 251178 472046 251274 472102
rect 251330 472046 251398 472102
rect 251454 472046 251522 472102
rect 251578 472046 251646 472102
rect 251702 472046 251798 472102
rect 251178 471978 251798 472046
rect 251178 471922 251274 471978
rect 251330 471922 251398 471978
rect 251454 471922 251522 471978
rect 251578 471922 251646 471978
rect 251702 471922 251798 471978
rect 251178 454350 251798 471922
rect 251178 454294 251274 454350
rect 251330 454294 251398 454350
rect 251454 454294 251522 454350
rect 251578 454294 251646 454350
rect 251702 454294 251798 454350
rect 251178 454226 251798 454294
rect 251178 454170 251274 454226
rect 251330 454170 251398 454226
rect 251454 454170 251522 454226
rect 251578 454170 251646 454226
rect 251702 454170 251798 454226
rect 251178 454102 251798 454170
rect 251178 454046 251274 454102
rect 251330 454046 251398 454102
rect 251454 454046 251522 454102
rect 251578 454046 251646 454102
rect 251702 454046 251798 454102
rect 251178 453978 251798 454046
rect 251178 453922 251274 453978
rect 251330 453922 251398 453978
rect 251454 453922 251522 453978
rect 251578 453922 251646 453978
rect 251702 453922 251798 453978
rect 251178 436350 251798 453922
rect 251178 436294 251274 436350
rect 251330 436294 251398 436350
rect 251454 436294 251522 436350
rect 251578 436294 251646 436350
rect 251702 436294 251798 436350
rect 251178 436226 251798 436294
rect 251178 436170 251274 436226
rect 251330 436170 251398 436226
rect 251454 436170 251522 436226
rect 251578 436170 251646 436226
rect 251702 436170 251798 436226
rect 251178 436102 251798 436170
rect 251178 436046 251274 436102
rect 251330 436046 251398 436102
rect 251454 436046 251522 436102
rect 251578 436046 251646 436102
rect 251702 436046 251798 436102
rect 251178 435978 251798 436046
rect 251178 435922 251274 435978
rect 251330 435922 251398 435978
rect 251454 435922 251522 435978
rect 251578 435922 251646 435978
rect 251702 435922 251798 435978
rect 249564 429268 249620 429278
rect 249564 427700 249620 429212
rect 249564 427634 249620 427644
rect 251178 425262 251798 435922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 568350 255518 585922
rect 254898 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 255518 568350
rect 254898 568226 255518 568294
rect 254898 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 255518 568226
rect 254898 568102 255518 568170
rect 254898 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 255518 568102
rect 254898 567978 255518 568046
rect 254898 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 255518 567978
rect 254898 550350 255518 567922
rect 254898 550294 254994 550350
rect 255050 550294 255118 550350
rect 255174 550294 255242 550350
rect 255298 550294 255366 550350
rect 255422 550294 255518 550350
rect 254898 550226 255518 550294
rect 254898 550170 254994 550226
rect 255050 550170 255118 550226
rect 255174 550170 255242 550226
rect 255298 550170 255366 550226
rect 255422 550170 255518 550226
rect 254898 550102 255518 550170
rect 254898 550046 254994 550102
rect 255050 550046 255118 550102
rect 255174 550046 255242 550102
rect 255298 550046 255366 550102
rect 255422 550046 255518 550102
rect 254898 549978 255518 550046
rect 254898 549922 254994 549978
rect 255050 549922 255118 549978
rect 255174 549922 255242 549978
rect 255298 549922 255366 549978
rect 255422 549922 255518 549978
rect 254898 532350 255518 549922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 281898 562350 282518 579922
rect 281898 562294 281994 562350
rect 282050 562294 282118 562350
rect 282174 562294 282242 562350
rect 282298 562294 282366 562350
rect 282422 562294 282518 562350
rect 281898 562226 282518 562294
rect 281898 562170 281994 562226
rect 282050 562170 282118 562226
rect 282174 562170 282242 562226
rect 282298 562170 282366 562226
rect 282422 562170 282518 562226
rect 281898 562102 282518 562170
rect 281898 562046 281994 562102
rect 282050 562046 282118 562102
rect 282174 562046 282242 562102
rect 282298 562046 282366 562102
rect 282422 562046 282518 562102
rect 281898 561978 282518 562046
rect 281898 561922 281994 561978
rect 282050 561922 282118 561978
rect 282174 561922 282242 561978
rect 282298 561922 282366 561978
rect 282422 561922 282518 561978
rect 268716 546418 268772 546428
rect 254898 532294 254994 532350
rect 255050 532294 255118 532350
rect 255174 532294 255242 532350
rect 255298 532294 255366 532350
rect 255422 532294 255518 532350
rect 254898 532226 255518 532294
rect 254898 532170 254994 532226
rect 255050 532170 255118 532226
rect 255174 532170 255242 532226
rect 255298 532170 255366 532226
rect 255422 532170 255518 532226
rect 254898 532102 255518 532170
rect 254898 532046 254994 532102
rect 255050 532046 255118 532102
rect 255174 532046 255242 532102
rect 255298 532046 255366 532102
rect 255422 532046 255518 532102
rect 254898 531978 255518 532046
rect 254898 531922 254994 531978
rect 255050 531922 255118 531978
rect 255174 531922 255242 531978
rect 255298 531922 255366 531978
rect 255422 531922 255518 531978
rect 254898 514350 255518 531922
rect 254898 514294 254994 514350
rect 255050 514294 255118 514350
rect 255174 514294 255242 514350
rect 255298 514294 255366 514350
rect 255422 514294 255518 514350
rect 254898 514226 255518 514294
rect 254898 514170 254994 514226
rect 255050 514170 255118 514226
rect 255174 514170 255242 514226
rect 255298 514170 255366 514226
rect 255422 514170 255518 514226
rect 254898 514102 255518 514170
rect 254898 514046 254994 514102
rect 255050 514046 255118 514102
rect 255174 514046 255242 514102
rect 255298 514046 255366 514102
rect 255422 514046 255518 514102
rect 254898 513978 255518 514046
rect 254898 513922 254994 513978
rect 255050 513922 255118 513978
rect 255174 513922 255242 513978
rect 255298 513922 255366 513978
rect 255422 513922 255518 513978
rect 254898 496350 255518 513922
rect 254898 496294 254994 496350
rect 255050 496294 255118 496350
rect 255174 496294 255242 496350
rect 255298 496294 255366 496350
rect 255422 496294 255518 496350
rect 254898 496226 255518 496294
rect 254898 496170 254994 496226
rect 255050 496170 255118 496226
rect 255174 496170 255242 496226
rect 255298 496170 255366 496226
rect 255422 496170 255518 496226
rect 254898 496102 255518 496170
rect 254898 496046 254994 496102
rect 255050 496046 255118 496102
rect 255174 496046 255242 496102
rect 255298 496046 255366 496102
rect 255422 496046 255518 496102
rect 254898 495978 255518 496046
rect 254898 495922 254994 495978
rect 255050 495922 255118 495978
rect 255174 495922 255242 495978
rect 255298 495922 255366 495978
rect 255422 495922 255518 495978
rect 254898 478350 255518 495922
rect 254898 478294 254994 478350
rect 255050 478294 255118 478350
rect 255174 478294 255242 478350
rect 255298 478294 255366 478350
rect 255422 478294 255518 478350
rect 254898 478226 255518 478294
rect 254898 478170 254994 478226
rect 255050 478170 255118 478226
rect 255174 478170 255242 478226
rect 255298 478170 255366 478226
rect 255422 478170 255518 478226
rect 254898 478102 255518 478170
rect 254898 478046 254994 478102
rect 255050 478046 255118 478102
rect 255174 478046 255242 478102
rect 255298 478046 255366 478102
rect 255422 478046 255518 478102
rect 254898 477978 255518 478046
rect 254898 477922 254994 477978
rect 255050 477922 255118 477978
rect 255174 477922 255242 477978
rect 255298 477922 255366 477978
rect 255422 477922 255518 477978
rect 254898 460350 255518 477922
rect 254898 460294 254994 460350
rect 255050 460294 255118 460350
rect 255174 460294 255242 460350
rect 255298 460294 255366 460350
rect 255422 460294 255518 460350
rect 254898 460226 255518 460294
rect 254898 460170 254994 460226
rect 255050 460170 255118 460226
rect 255174 460170 255242 460226
rect 255298 460170 255366 460226
rect 255422 460170 255518 460226
rect 254898 460102 255518 460170
rect 254898 460046 254994 460102
rect 255050 460046 255118 460102
rect 255174 460046 255242 460102
rect 255298 460046 255366 460102
rect 255422 460046 255518 460102
rect 254898 459978 255518 460046
rect 254898 459922 254994 459978
rect 255050 459922 255118 459978
rect 255174 459922 255242 459978
rect 255298 459922 255366 459978
rect 255422 459922 255518 459978
rect 254898 442350 255518 459922
rect 254898 442294 254994 442350
rect 255050 442294 255118 442350
rect 255174 442294 255242 442350
rect 255298 442294 255366 442350
rect 255422 442294 255518 442350
rect 254898 442226 255518 442294
rect 254898 442170 254994 442226
rect 255050 442170 255118 442226
rect 255174 442170 255242 442226
rect 255298 442170 255366 442226
rect 255422 442170 255518 442226
rect 254898 442102 255518 442170
rect 254898 442046 254994 442102
rect 255050 442046 255118 442102
rect 255174 442046 255242 442102
rect 255298 442046 255366 442102
rect 255422 442046 255518 442102
rect 254898 441978 255518 442046
rect 254898 441922 254994 441978
rect 255050 441922 255118 441978
rect 255174 441922 255242 441978
rect 255298 441922 255366 441978
rect 255422 441922 255518 441978
rect 252252 429268 252308 429278
rect 252252 427812 252308 429212
rect 252252 427746 252308 427756
rect 254898 425262 255518 441922
rect 267036 546238 267092 546248
rect 267036 433412 267092 546182
rect 267036 433346 267092 433356
rect 268716 433412 268772 546362
rect 268716 433346 268772 433356
rect 281898 544350 282518 561922
rect 281898 544294 281994 544350
rect 282050 544294 282118 544350
rect 282174 544294 282242 544350
rect 282298 544294 282366 544350
rect 282422 544294 282518 544350
rect 281898 544226 282518 544294
rect 281898 544170 281994 544226
rect 282050 544170 282118 544226
rect 282174 544170 282242 544226
rect 282298 544170 282366 544226
rect 282422 544170 282518 544226
rect 281898 544102 282518 544170
rect 281898 544046 281994 544102
rect 282050 544046 282118 544102
rect 282174 544046 282242 544102
rect 282298 544046 282366 544102
rect 282422 544046 282518 544102
rect 281898 543978 282518 544046
rect 281898 543922 281994 543978
rect 282050 543922 282118 543978
rect 282174 543922 282242 543978
rect 282298 543922 282366 543978
rect 282422 543922 282518 543978
rect 281898 526350 282518 543922
rect 281898 526294 281994 526350
rect 282050 526294 282118 526350
rect 282174 526294 282242 526350
rect 282298 526294 282366 526350
rect 282422 526294 282518 526350
rect 281898 526226 282518 526294
rect 281898 526170 281994 526226
rect 282050 526170 282118 526226
rect 282174 526170 282242 526226
rect 282298 526170 282366 526226
rect 282422 526170 282518 526226
rect 281898 526102 282518 526170
rect 281898 526046 281994 526102
rect 282050 526046 282118 526102
rect 282174 526046 282242 526102
rect 282298 526046 282366 526102
rect 282422 526046 282518 526102
rect 281898 525978 282518 526046
rect 281898 525922 281994 525978
rect 282050 525922 282118 525978
rect 282174 525922 282242 525978
rect 282298 525922 282366 525978
rect 282422 525922 282518 525978
rect 281898 508350 282518 525922
rect 281898 508294 281994 508350
rect 282050 508294 282118 508350
rect 282174 508294 282242 508350
rect 282298 508294 282366 508350
rect 282422 508294 282518 508350
rect 281898 508226 282518 508294
rect 281898 508170 281994 508226
rect 282050 508170 282118 508226
rect 282174 508170 282242 508226
rect 282298 508170 282366 508226
rect 282422 508170 282518 508226
rect 281898 508102 282518 508170
rect 281898 508046 281994 508102
rect 282050 508046 282118 508102
rect 282174 508046 282242 508102
rect 282298 508046 282366 508102
rect 282422 508046 282518 508102
rect 281898 507978 282518 508046
rect 281898 507922 281994 507978
rect 282050 507922 282118 507978
rect 282174 507922 282242 507978
rect 282298 507922 282366 507978
rect 282422 507922 282518 507978
rect 281898 490350 282518 507922
rect 281898 490294 281994 490350
rect 282050 490294 282118 490350
rect 282174 490294 282242 490350
rect 282298 490294 282366 490350
rect 282422 490294 282518 490350
rect 281898 490226 282518 490294
rect 281898 490170 281994 490226
rect 282050 490170 282118 490226
rect 282174 490170 282242 490226
rect 282298 490170 282366 490226
rect 282422 490170 282518 490226
rect 281898 490102 282518 490170
rect 281898 490046 281994 490102
rect 282050 490046 282118 490102
rect 282174 490046 282242 490102
rect 282298 490046 282366 490102
rect 282422 490046 282518 490102
rect 281898 489978 282518 490046
rect 281898 489922 281994 489978
rect 282050 489922 282118 489978
rect 282174 489922 282242 489978
rect 282298 489922 282366 489978
rect 282422 489922 282518 489978
rect 281898 472350 282518 489922
rect 281898 472294 281994 472350
rect 282050 472294 282118 472350
rect 282174 472294 282242 472350
rect 282298 472294 282366 472350
rect 282422 472294 282518 472350
rect 281898 472226 282518 472294
rect 281898 472170 281994 472226
rect 282050 472170 282118 472226
rect 282174 472170 282242 472226
rect 282298 472170 282366 472226
rect 282422 472170 282518 472226
rect 281898 472102 282518 472170
rect 281898 472046 281994 472102
rect 282050 472046 282118 472102
rect 282174 472046 282242 472102
rect 282298 472046 282366 472102
rect 282422 472046 282518 472102
rect 281898 471978 282518 472046
rect 281898 471922 281994 471978
rect 282050 471922 282118 471978
rect 282174 471922 282242 471978
rect 282298 471922 282366 471978
rect 282422 471922 282518 471978
rect 281898 454350 282518 471922
rect 281898 454294 281994 454350
rect 282050 454294 282118 454350
rect 282174 454294 282242 454350
rect 282298 454294 282366 454350
rect 282422 454294 282518 454350
rect 281898 454226 282518 454294
rect 281898 454170 281994 454226
rect 282050 454170 282118 454226
rect 282174 454170 282242 454226
rect 282298 454170 282366 454226
rect 282422 454170 282518 454226
rect 281898 454102 282518 454170
rect 281898 454046 281994 454102
rect 282050 454046 282118 454102
rect 282174 454046 282242 454102
rect 282298 454046 282366 454102
rect 282422 454046 282518 454102
rect 281898 453978 282518 454046
rect 281898 453922 281994 453978
rect 282050 453922 282118 453978
rect 282174 453922 282242 453978
rect 282298 453922 282366 453978
rect 282422 453922 282518 453978
rect 281898 436350 282518 453922
rect 281898 436294 281994 436350
rect 282050 436294 282118 436350
rect 282174 436294 282242 436350
rect 282298 436294 282366 436350
rect 282422 436294 282518 436350
rect 281898 436226 282518 436294
rect 281898 436170 281994 436226
rect 282050 436170 282118 436226
rect 282174 436170 282242 436226
rect 282298 436170 282366 436226
rect 282422 436170 282518 436226
rect 281898 436102 282518 436170
rect 281898 436046 281994 436102
rect 282050 436046 282118 436102
rect 282174 436046 282242 436102
rect 282298 436046 282366 436102
rect 282422 436046 282518 436102
rect 281898 435978 282518 436046
rect 281898 435922 281994 435978
rect 282050 435922 282118 435978
rect 282174 435922 282242 435978
rect 282298 435922 282366 435978
rect 282422 435922 282518 435978
rect 276332 432118 276388 432128
rect 260316 429268 260372 429278
rect 110528 424350 110848 424384
rect 110528 424294 110598 424350
rect 110654 424294 110722 424350
rect 110778 424294 110848 424350
rect 110528 424226 110848 424294
rect 110528 424170 110598 424226
rect 110654 424170 110722 424226
rect 110778 424170 110848 424226
rect 110528 424102 110848 424170
rect 110528 424046 110598 424102
rect 110654 424046 110722 424102
rect 110778 424046 110848 424102
rect 110528 423978 110848 424046
rect 110528 423922 110598 423978
rect 110654 423922 110722 423978
rect 110778 423922 110848 423978
rect 110528 423888 110848 423922
rect 141248 424350 141568 424384
rect 141248 424294 141318 424350
rect 141374 424294 141442 424350
rect 141498 424294 141568 424350
rect 141248 424226 141568 424294
rect 141248 424170 141318 424226
rect 141374 424170 141442 424226
rect 141498 424170 141568 424226
rect 141248 424102 141568 424170
rect 141248 424046 141318 424102
rect 141374 424046 141442 424102
rect 141498 424046 141568 424102
rect 141248 423978 141568 424046
rect 141248 423922 141318 423978
rect 141374 423922 141442 423978
rect 141498 423922 141568 423978
rect 141248 423888 141568 423922
rect 171968 424350 172288 424384
rect 171968 424294 172038 424350
rect 172094 424294 172162 424350
rect 172218 424294 172288 424350
rect 171968 424226 172288 424294
rect 171968 424170 172038 424226
rect 172094 424170 172162 424226
rect 172218 424170 172288 424226
rect 171968 424102 172288 424170
rect 171968 424046 172038 424102
rect 172094 424046 172162 424102
rect 172218 424046 172288 424102
rect 171968 423978 172288 424046
rect 171968 423922 172038 423978
rect 172094 423922 172162 423978
rect 172218 423922 172288 423978
rect 171968 423888 172288 423922
rect 202688 424350 203008 424384
rect 202688 424294 202758 424350
rect 202814 424294 202882 424350
rect 202938 424294 203008 424350
rect 202688 424226 203008 424294
rect 202688 424170 202758 424226
rect 202814 424170 202882 424226
rect 202938 424170 203008 424226
rect 202688 424102 203008 424170
rect 202688 424046 202758 424102
rect 202814 424046 202882 424102
rect 202938 424046 203008 424102
rect 202688 423978 203008 424046
rect 202688 423922 202758 423978
rect 202814 423922 202882 423978
rect 202938 423922 203008 423978
rect 202688 423888 203008 423922
rect 233408 424350 233728 424384
rect 233408 424294 233478 424350
rect 233534 424294 233602 424350
rect 233658 424294 233728 424350
rect 233408 424226 233728 424294
rect 233408 424170 233478 424226
rect 233534 424170 233602 424226
rect 233658 424170 233728 424226
rect 233408 424102 233728 424170
rect 233408 424046 233478 424102
rect 233534 424046 233602 424102
rect 233658 424046 233728 424102
rect 233408 423978 233728 424046
rect 233408 423922 233478 423978
rect 233534 423922 233602 423978
rect 233658 423922 233728 423978
rect 233408 423888 233728 423922
rect 95168 418350 95488 418384
rect 95168 418294 95238 418350
rect 95294 418294 95362 418350
rect 95418 418294 95488 418350
rect 95168 418226 95488 418294
rect 95168 418170 95238 418226
rect 95294 418170 95362 418226
rect 95418 418170 95488 418226
rect 95168 418102 95488 418170
rect 95168 418046 95238 418102
rect 95294 418046 95362 418102
rect 95418 418046 95488 418102
rect 95168 417978 95488 418046
rect 95168 417922 95238 417978
rect 95294 417922 95362 417978
rect 95418 417922 95488 417978
rect 95168 417888 95488 417922
rect 125888 418350 126208 418384
rect 125888 418294 125958 418350
rect 126014 418294 126082 418350
rect 126138 418294 126208 418350
rect 125888 418226 126208 418294
rect 125888 418170 125958 418226
rect 126014 418170 126082 418226
rect 126138 418170 126208 418226
rect 125888 418102 126208 418170
rect 125888 418046 125958 418102
rect 126014 418046 126082 418102
rect 126138 418046 126208 418102
rect 125888 417978 126208 418046
rect 125888 417922 125958 417978
rect 126014 417922 126082 417978
rect 126138 417922 126208 417978
rect 125888 417888 126208 417922
rect 156608 418350 156928 418384
rect 156608 418294 156678 418350
rect 156734 418294 156802 418350
rect 156858 418294 156928 418350
rect 156608 418226 156928 418294
rect 156608 418170 156678 418226
rect 156734 418170 156802 418226
rect 156858 418170 156928 418226
rect 156608 418102 156928 418170
rect 156608 418046 156678 418102
rect 156734 418046 156802 418102
rect 156858 418046 156928 418102
rect 156608 417978 156928 418046
rect 156608 417922 156678 417978
rect 156734 417922 156802 417978
rect 156858 417922 156928 417978
rect 156608 417888 156928 417922
rect 187328 418350 187648 418384
rect 187328 418294 187398 418350
rect 187454 418294 187522 418350
rect 187578 418294 187648 418350
rect 187328 418226 187648 418294
rect 187328 418170 187398 418226
rect 187454 418170 187522 418226
rect 187578 418170 187648 418226
rect 187328 418102 187648 418170
rect 187328 418046 187398 418102
rect 187454 418046 187522 418102
rect 187578 418046 187648 418102
rect 187328 417978 187648 418046
rect 187328 417922 187398 417978
rect 187454 417922 187522 417978
rect 187578 417922 187648 417978
rect 187328 417888 187648 417922
rect 218048 418350 218368 418384
rect 218048 418294 218118 418350
rect 218174 418294 218242 418350
rect 218298 418294 218368 418350
rect 218048 418226 218368 418294
rect 218048 418170 218118 418226
rect 218174 418170 218242 418226
rect 218298 418170 218368 418226
rect 218048 418102 218368 418170
rect 218048 418046 218118 418102
rect 218174 418046 218242 418102
rect 218298 418046 218368 418102
rect 218048 417978 218368 418046
rect 218048 417922 218118 417978
rect 218174 417922 218242 417978
rect 218298 417922 218368 417978
rect 218048 417888 218368 417922
rect 248768 418350 249088 418384
rect 248768 418294 248838 418350
rect 248894 418294 248962 418350
rect 249018 418294 249088 418350
rect 248768 418226 249088 418294
rect 248768 418170 248838 418226
rect 248894 418170 248962 418226
rect 249018 418170 249088 418226
rect 248768 418102 249088 418170
rect 248768 418046 248838 418102
rect 248894 418046 248962 418102
rect 249018 418046 249088 418102
rect 248768 417978 249088 418046
rect 248768 417922 248838 417978
rect 248894 417922 248962 417978
rect 249018 417922 249088 417978
rect 248768 417888 249088 417922
rect 83580 409732 83636 409742
rect 110528 406350 110848 406384
rect 110528 406294 110598 406350
rect 110654 406294 110722 406350
rect 110778 406294 110848 406350
rect 110528 406226 110848 406294
rect 110528 406170 110598 406226
rect 110654 406170 110722 406226
rect 110778 406170 110848 406226
rect 110528 406102 110848 406170
rect 110528 406046 110598 406102
rect 110654 406046 110722 406102
rect 110778 406046 110848 406102
rect 110528 405978 110848 406046
rect 110528 405922 110598 405978
rect 110654 405922 110722 405978
rect 110778 405922 110848 405978
rect 110528 405888 110848 405922
rect 141248 406350 141568 406384
rect 141248 406294 141318 406350
rect 141374 406294 141442 406350
rect 141498 406294 141568 406350
rect 141248 406226 141568 406294
rect 141248 406170 141318 406226
rect 141374 406170 141442 406226
rect 141498 406170 141568 406226
rect 141248 406102 141568 406170
rect 141248 406046 141318 406102
rect 141374 406046 141442 406102
rect 141498 406046 141568 406102
rect 141248 405978 141568 406046
rect 141248 405922 141318 405978
rect 141374 405922 141442 405978
rect 141498 405922 141568 405978
rect 141248 405888 141568 405922
rect 171968 406350 172288 406384
rect 171968 406294 172038 406350
rect 172094 406294 172162 406350
rect 172218 406294 172288 406350
rect 171968 406226 172288 406294
rect 171968 406170 172038 406226
rect 172094 406170 172162 406226
rect 172218 406170 172288 406226
rect 171968 406102 172288 406170
rect 171968 406046 172038 406102
rect 172094 406046 172162 406102
rect 172218 406046 172288 406102
rect 171968 405978 172288 406046
rect 171968 405922 172038 405978
rect 172094 405922 172162 405978
rect 172218 405922 172288 405978
rect 171968 405888 172288 405922
rect 202688 406350 203008 406384
rect 202688 406294 202758 406350
rect 202814 406294 202882 406350
rect 202938 406294 203008 406350
rect 202688 406226 203008 406294
rect 202688 406170 202758 406226
rect 202814 406170 202882 406226
rect 202938 406170 203008 406226
rect 202688 406102 203008 406170
rect 202688 406046 202758 406102
rect 202814 406046 202882 406102
rect 202938 406046 203008 406102
rect 202688 405978 203008 406046
rect 202688 405922 202758 405978
rect 202814 405922 202882 405978
rect 202938 405922 203008 405978
rect 202688 405888 203008 405922
rect 233408 406350 233728 406384
rect 233408 406294 233478 406350
rect 233534 406294 233602 406350
rect 233658 406294 233728 406350
rect 233408 406226 233728 406294
rect 233408 406170 233478 406226
rect 233534 406170 233602 406226
rect 233658 406170 233728 406226
rect 233408 406102 233728 406170
rect 233408 406046 233478 406102
rect 233534 406046 233602 406102
rect 233658 406046 233728 406102
rect 233408 405978 233728 406046
rect 233408 405922 233478 405978
rect 233534 405922 233602 405978
rect 233658 405922 233728 405978
rect 233408 405888 233728 405922
rect 260316 403138 260372 429212
rect 260316 403072 260372 403082
rect 263676 429268 263732 429278
rect 263676 402958 263732 429212
rect 264128 424350 264448 424384
rect 264128 424294 264198 424350
rect 264254 424294 264322 424350
rect 264378 424294 264448 424350
rect 264128 424226 264448 424294
rect 264128 424170 264198 424226
rect 264254 424170 264322 424226
rect 264378 424170 264448 424226
rect 264128 424102 264448 424170
rect 264128 424046 264198 424102
rect 264254 424046 264322 424102
rect 264378 424046 264448 424102
rect 264128 423978 264448 424046
rect 264128 423922 264198 423978
rect 264254 423922 264322 423978
rect 264378 423922 264448 423978
rect 264128 423888 264448 423922
rect 264128 406350 264448 406384
rect 264128 406294 264198 406350
rect 264254 406294 264322 406350
rect 264378 406294 264448 406350
rect 264128 406226 264448 406294
rect 264128 406170 264198 406226
rect 264254 406170 264322 406226
rect 264378 406170 264448 406226
rect 264128 406102 264448 406170
rect 264128 406046 264198 406102
rect 264254 406046 264322 406102
rect 264378 406046 264448 406102
rect 264128 405978 264448 406046
rect 264128 405922 264198 405978
rect 264254 405922 264322 405978
rect 264378 405922 264448 405978
rect 264128 405888 264448 405922
rect 263676 402892 263732 402902
rect 95168 400350 95488 400384
rect 95168 400294 95238 400350
rect 95294 400294 95362 400350
rect 95418 400294 95488 400350
rect 95168 400226 95488 400294
rect 95168 400170 95238 400226
rect 95294 400170 95362 400226
rect 95418 400170 95488 400226
rect 95168 400102 95488 400170
rect 95168 400046 95238 400102
rect 95294 400046 95362 400102
rect 95418 400046 95488 400102
rect 95168 399978 95488 400046
rect 95168 399922 95238 399978
rect 95294 399922 95362 399978
rect 95418 399922 95488 399978
rect 95168 399888 95488 399922
rect 125888 400350 126208 400384
rect 125888 400294 125958 400350
rect 126014 400294 126082 400350
rect 126138 400294 126208 400350
rect 125888 400226 126208 400294
rect 125888 400170 125958 400226
rect 126014 400170 126082 400226
rect 126138 400170 126208 400226
rect 125888 400102 126208 400170
rect 125888 400046 125958 400102
rect 126014 400046 126082 400102
rect 126138 400046 126208 400102
rect 125888 399978 126208 400046
rect 125888 399922 125958 399978
rect 126014 399922 126082 399978
rect 126138 399922 126208 399978
rect 125888 399888 126208 399922
rect 156608 400350 156928 400384
rect 156608 400294 156678 400350
rect 156734 400294 156802 400350
rect 156858 400294 156928 400350
rect 156608 400226 156928 400294
rect 156608 400170 156678 400226
rect 156734 400170 156802 400226
rect 156858 400170 156928 400226
rect 156608 400102 156928 400170
rect 156608 400046 156678 400102
rect 156734 400046 156802 400102
rect 156858 400046 156928 400102
rect 156608 399978 156928 400046
rect 156608 399922 156678 399978
rect 156734 399922 156802 399978
rect 156858 399922 156928 399978
rect 156608 399888 156928 399922
rect 187328 400350 187648 400384
rect 187328 400294 187398 400350
rect 187454 400294 187522 400350
rect 187578 400294 187648 400350
rect 187328 400226 187648 400294
rect 187328 400170 187398 400226
rect 187454 400170 187522 400226
rect 187578 400170 187648 400226
rect 187328 400102 187648 400170
rect 187328 400046 187398 400102
rect 187454 400046 187522 400102
rect 187578 400046 187648 400102
rect 187328 399978 187648 400046
rect 187328 399922 187398 399978
rect 187454 399922 187522 399978
rect 187578 399922 187648 399978
rect 187328 399888 187648 399922
rect 218048 400350 218368 400384
rect 218048 400294 218118 400350
rect 218174 400294 218242 400350
rect 218298 400294 218368 400350
rect 218048 400226 218368 400294
rect 218048 400170 218118 400226
rect 218174 400170 218242 400226
rect 218298 400170 218368 400226
rect 218048 400102 218368 400170
rect 218048 400046 218118 400102
rect 218174 400046 218242 400102
rect 218298 400046 218368 400102
rect 218048 399978 218368 400046
rect 218048 399922 218118 399978
rect 218174 399922 218242 399978
rect 218298 399922 218368 399978
rect 218048 399888 218368 399922
rect 248768 400350 249088 400384
rect 248768 400294 248838 400350
rect 248894 400294 248962 400350
rect 249018 400294 249088 400350
rect 248768 400226 249088 400294
rect 248768 400170 248838 400226
rect 248894 400170 248962 400226
rect 249018 400170 249088 400226
rect 248768 400102 249088 400170
rect 248768 400046 248838 400102
rect 248894 400046 248962 400102
rect 249018 400046 249088 400102
rect 248768 399978 249088 400046
rect 248768 399922 248838 399978
rect 248894 399922 248962 399978
rect 249018 399922 249088 399978
rect 248768 399888 249088 399922
rect 273196 390628 273252 390638
rect 110528 388350 110848 388384
rect 110528 388294 110598 388350
rect 110654 388294 110722 388350
rect 110778 388294 110848 388350
rect 110528 388226 110848 388294
rect 110528 388170 110598 388226
rect 110654 388170 110722 388226
rect 110778 388170 110848 388226
rect 110528 388102 110848 388170
rect 110528 388046 110598 388102
rect 110654 388046 110722 388102
rect 110778 388046 110848 388102
rect 110528 387978 110848 388046
rect 110528 387922 110598 387978
rect 110654 387922 110722 387978
rect 110778 387922 110848 387978
rect 110528 387888 110848 387922
rect 141248 388350 141568 388384
rect 141248 388294 141318 388350
rect 141374 388294 141442 388350
rect 141498 388294 141568 388350
rect 141248 388226 141568 388294
rect 141248 388170 141318 388226
rect 141374 388170 141442 388226
rect 141498 388170 141568 388226
rect 141248 388102 141568 388170
rect 141248 388046 141318 388102
rect 141374 388046 141442 388102
rect 141498 388046 141568 388102
rect 141248 387978 141568 388046
rect 141248 387922 141318 387978
rect 141374 387922 141442 387978
rect 141498 387922 141568 387978
rect 141248 387888 141568 387922
rect 171968 388350 172288 388384
rect 171968 388294 172038 388350
rect 172094 388294 172162 388350
rect 172218 388294 172288 388350
rect 171968 388226 172288 388294
rect 171968 388170 172038 388226
rect 172094 388170 172162 388226
rect 172218 388170 172288 388226
rect 171968 388102 172288 388170
rect 171968 388046 172038 388102
rect 172094 388046 172162 388102
rect 172218 388046 172288 388102
rect 171968 387978 172288 388046
rect 171968 387922 172038 387978
rect 172094 387922 172162 387978
rect 172218 387922 172288 387978
rect 171968 387888 172288 387922
rect 202688 388350 203008 388384
rect 202688 388294 202758 388350
rect 202814 388294 202882 388350
rect 202938 388294 203008 388350
rect 202688 388226 203008 388294
rect 202688 388170 202758 388226
rect 202814 388170 202882 388226
rect 202938 388170 203008 388226
rect 202688 388102 203008 388170
rect 202688 388046 202758 388102
rect 202814 388046 202882 388102
rect 202938 388046 203008 388102
rect 202688 387978 203008 388046
rect 202688 387922 202758 387978
rect 202814 387922 202882 387978
rect 202938 387922 203008 387978
rect 202688 387888 203008 387922
rect 233408 388350 233728 388384
rect 233408 388294 233478 388350
rect 233534 388294 233602 388350
rect 233658 388294 233728 388350
rect 233408 388226 233728 388294
rect 233408 388170 233478 388226
rect 233534 388170 233602 388226
rect 233658 388170 233728 388226
rect 233408 388102 233728 388170
rect 233408 388046 233478 388102
rect 233534 388046 233602 388102
rect 233658 388046 233728 388102
rect 233408 387978 233728 388046
rect 233408 387922 233478 387978
rect 233534 387922 233602 387978
rect 233658 387922 233728 387978
rect 233408 387888 233728 387922
rect 264128 388350 264448 388384
rect 264128 388294 264198 388350
rect 264254 388294 264322 388350
rect 264378 388294 264448 388350
rect 264128 388226 264448 388294
rect 264128 388170 264198 388226
rect 264254 388170 264322 388226
rect 264378 388170 264448 388226
rect 264128 388102 264448 388170
rect 264128 388046 264198 388102
rect 264254 388046 264322 388102
rect 264378 388046 264448 388102
rect 264128 387978 264448 388046
rect 264128 387922 264198 387978
rect 264254 387922 264322 387978
rect 264378 387922 264448 387978
rect 264128 387888 264448 387922
rect 84812 383158 84868 383168
rect 83468 347632 83524 347642
rect 83580 368218 83636 368228
rect 83580 295318 83636 368162
rect 83804 368038 83860 368048
rect 83580 295252 83636 295262
rect 83692 366418 83748 366428
rect 83692 295138 83748 366362
rect 83804 298918 83860 367982
rect 84812 300178 84868 383102
rect 95168 382350 95488 382384
rect 95168 382294 95238 382350
rect 95294 382294 95362 382350
rect 95418 382294 95488 382350
rect 95168 382226 95488 382294
rect 95168 382170 95238 382226
rect 95294 382170 95362 382226
rect 95418 382170 95488 382226
rect 95168 382102 95488 382170
rect 95168 382046 95238 382102
rect 95294 382046 95362 382102
rect 95418 382046 95488 382102
rect 95168 381978 95488 382046
rect 95168 381922 95238 381978
rect 95294 381922 95362 381978
rect 95418 381922 95488 381978
rect 95168 381888 95488 381922
rect 125888 382350 126208 382384
rect 125888 382294 125958 382350
rect 126014 382294 126082 382350
rect 126138 382294 126208 382350
rect 125888 382226 126208 382294
rect 125888 382170 125958 382226
rect 126014 382170 126082 382226
rect 126138 382170 126208 382226
rect 125888 382102 126208 382170
rect 125888 382046 125958 382102
rect 126014 382046 126082 382102
rect 126138 382046 126208 382102
rect 125888 381978 126208 382046
rect 125888 381922 125958 381978
rect 126014 381922 126082 381978
rect 126138 381922 126208 381978
rect 125888 381888 126208 381922
rect 156608 382350 156928 382384
rect 156608 382294 156678 382350
rect 156734 382294 156802 382350
rect 156858 382294 156928 382350
rect 156608 382226 156928 382294
rect 156608 382170 156678 382226
rect 156734 382170 156802 382226
rect 156858 382170 156928 382226
rect 156608 382102 156928 382170
rect 156608 382046 156678 382102
rect 156734 382046 156802 382102
rect 156858 382046 156928 382102
rect 156608 381978 156928 382046
rect 156608 381922 156678 381978
rect 156734 381922 156802 381978
rect 156858 381922 156928 381978
rect 156608 381888 156928 381922
rect 187328 382350 187648 382384
rect 187328 382294 187398 382350
rect 187454 382294 187522 382350
rect 187578 382294 187648 382350
rect 187328 382226 187648 382294
rect 187328 382170 187398 382226
rect 187454 382170 187522 382226
rect 187578 382170 187648 382226
rect 187328 382102 187648 382170
rect 187328 382046 187398 382102
rect 187454 382046 187522 382102
rect 187578 382046 187648 382102
rect 187328 381978 187648 382046
rect 187328 381922 187398 381978
rect 187454 381922 187522 381978
rect 187578 381922 187648 381978
rect 187328 381888 187648 381922
rect 218048 382350 218368 382384
rect 218048 382294 218118 382350
rect 218174 382294 218242 382350
rect 218298 382294 218368 382350
rect 218048 382226 218368 382294
rect 218048 382170 218118 382226
rect 218174 382170 218242 382226
rect 218298 382170 218368 382226
rect 218048 382102 218368 382170
rect 218048 382046 218118 382102
rect 218174 382046 218242 382102
rect 218298 382046 218368 382102
rect 218048 381978 218368 382046
rect 218048 381922 218118 381978
rect 218174 381922 218242 381978
rect 218298 381922 218368 381978
rect 218048 381888 218368 381922
rect 248768 382350 249088 382384
rect 248768 382294 248838 382350
rect 248894 382294 248962 382350
rect 249018 382294 249088 382350
rect 248768 382226 249088 382294
rect 248768 382170 248838 382226
rect 248894 382170 248962 382226
rect 249018 382170 249088 382226
rect 248768 382102 249088 382170
rect 248768 382046 248838 382102
rect 248894 382046 248962 382102
rect 249018 382046 249088 382102
rect 273196 382116 273252 390572
rect 273532 388918 273588 388928
rect 273532 388836 273588 388862
rect 273532 388770 273588 388780
rect 273196 382050 273252 382060
rect 273644 384020 273700 384030
rect 248768 381978 249088 382046
rect 248768 381922 248838 381978
rect 248894 381922 248962 381978
rect 249018 381922 249088 381978
rect 248768 381888 249088 381922
rect 273644 379428 273700 383964
rect 273644 379362 273700 379372
rect 273756 380660 273812 380670
rect 273756 378084 273812 380604
rect 276332 378868 276388 432062
rect 276444 432068 276500 432078
rect 276444 387658 276500 432012
rect 276444 387592 276500 387602
rect 278012 430612 278068 430622
rect 276332 378802 276388 378812
rect 273756 378018 273812 378028
rect 273756 371458 273812 371468
rect 273756 371364 273812 371402
rect 273756 371298 273812 371308
rect 110528 370350 110848 370384
rect 110528 370294 110598 370350
rect 110654 370294 110722 370350
rect 110778 370294 110848 370350
rect 110528 370226 110848 370294
rect 110528 370170 110598 370226
rect 110654 370170 110722 370226
rect 110778 370170 110848 370226
rect 110528 370102 110848 370170
rect 110528 370046 110598 370102
rect 110654 370046 110722 370102
rect 110778 370046 110848 370102
rect 110528 369978 110848 370046
rect 110528 369922 110598 369978
rect 110654 369922 110722 369978
rect 110778 369922 110848 369978
rect 110528 369888 110848 369922
rect 141248 370350 141568 370384
rect 141248 370294 141318 370350
rect 141374 370294 141442 370350
rect 141498 370294 141568 370350
rect 141248 370226 141568 370294
rect 141248 370170 141318 370226
rect 141374 370170 141442 370226
rect 141498 370170 141568 370226
rect 141248 370102 141568 370170
rect 141248 370046 141318 370102
rect 141374 370046 141442 370102
rect 141498 370046 141568 370102
rect 141248 369978 141568 370046
rect 141248 369922 141318 369978
rect 141374 369922 141442 369978
rect 141498 369922 141568 369978
rect 141248 369888 141568 369922
rect 171968 370350 172288 370384
rect 171968 370294 172038 370350
rect 172094 370294 172162 370350
rect 172218 370294 172288 370350
rect 171968 370226 172288 370294
rect 171968 370170 172038 370226
rect 172094 370170 172162 370226
rect 172218 370170 172288 370226
rect 171968 370102 172288 370170
rect 171968 370046 172038 370102
rect 172094 370046 172162 370102
rect 172218 370046 172288 370102
rect 171968 369978 172288 370046
rect 171968 369922 172038 369978
rect 172094 369922 172162 369978
rect 172218 369922 172288 369978
rect 171968 369888 172288 369922
rect 202688 370350 203008 370384
rect 202688 370294 202758 370350
rect 202814 370294 202882 370350
rect 202938 370294 203008 370350
rect 202688 370226 203008 370294
rect 202688 370170 202758 370226
rect 202814 370170 202882 370226
rect 202938 370170 203008 370226
rect 202688 370102 203008 370170
rect 202688 370046 202758 370102
rect 202814 370046 202882 370102
rect 202938 370046 203008 370102
rect 202688 369978 203008 370046
rect 202688 369922 202758 369978
rect 202814 369922 202882 369978
rect 202938 369922 203008 369978
rect 202688 369888 203008 369922
rect 233408 370350 233728 370384
rect 233408 370294 233478 370350
rect 233534 370294 233602 370350
rect 233658 370294 233728 370350
rect 233408 370226 233728 370294
rect 233408 370170 233478 370226
rect 233534 370170 233602 370226
rect 233658 370170 233728 370226
rect 233408 370102 233728 370170
rect 233408 370046 233478 370102
rect 233534 370046 233602 370102
rect 233658 370046 233728 370102
rect 233408 369978 233728 370046
rect 233408 369922 233478 369978
rect 233534 369922 233602 369978
rect 233658 369922 233728 369978
rect 233408 369888 233728 369922
rect 264128 370350 264448 370384
rect 264128 370294 264198 370350
rect 264254 370294 264322 370350
rect 264378 370294 264448 370350
rect 264128 370226 264448 370294
rect 264128 370170 264198 370226
rect 264254 370170 264322 370226
rect 264378 370170 264448 370226
rect 264128 370102 264448 370170
rect 264128 370046 264198 370102
rect 264254 370046 264322 370102
rect 264378 370046 264448 370102
rect 264128 369978 264448 370046
rect 264128 369922 264198 369978
rect 264254 369922 264322 369978
rect 264378 369922 264448 369978
rect 264128 369888 264448 369922
rect 273756 368676 273812 368686
rect 273756 368038 273812 368620
rect 273756 367972 273812 367982
rect 273756 367332 273812 367342
rect 273756 366418 273812 367276
rect 273756 366352 273812 366362
rect 273756 365988 273812 365998
rect 273756 364798 273812 365932
rect 273756 364732 273812 364742
rect 273756 364644 273812 364656
rect 273756 364552 273812 364562
rect 95168 364350 95488 364384
rect 95168 364294 95238 364350
rect 95294 364294 95362 364350
rect 95418 364294 95488 364350
rect 95168 364226 95488 364294
rect 95168 364170 95238 364226
rect 95294 364170 95362 364226
rect 95418 364170 95488 364226
rect 95168 364102 95488 364170
rect 95168 364046 95238 364102
rect 95294 364046 95362 364102
rect 95418 364046 95488 364102
rect 95168 363978 95488 364046
rect 95168 363922 95238 363978
rect 95294 363922 95362 363978
rect 95418 363922 95488 363978
rect 95168 363888 95488 363922
rect 125888 364350 126208 364384
rect 125888 364294 125958 364350
rect 126014 364294 126082 364350
rect 126138 364294 126208 364350
rect 125888 364226 126208 364294
rect 125888 364170 125958 364226
rect 126014 364170 126082 364226
rect 126138 364170 126208 364226
rect 125888 364102 126208 364170
rect 125888 364046 125958 364102
rect 126014 364046 126082 364102
rect 126138 364046 126208 364102
rect 125888 363978 126208 364046
rect 125888 363922 125958 363978
rect 126014 363922 126082 363978
rect 126138 363922 126208 363978
rect 125888 363888 126208 363922
rect 156608 364350 156928 364384
rect 156608 364294 156678 364350
rect 156734 364294 156802 364350
rect 156858 364294 156928 364350
rect 156608 364226 156928 364294
rect 156608 364170 156678 364226
rect 156734 364170 156802 364226
rect 156858 364170 156928 364226
rect 156608 364102 156928 364170
rect 156608 364046 156678 364102
rect 156734 364046 156802 364102
rect 156858 364046 156928 364102
rect 156608 363978 156928 364046
rect 156608 363922 156678 363978
rect 156734 363922 156802 363978
rect 156858 363922 156928 363978
rect 156608 363888 156928 363922
rect 187328 364350 187648 364384
rect 187328 364294 187398 364350
rect 187454 364294 187522 364350
rect 187578 364294 187648 364350
rect 187328 364226 187648 364294
rect 187328 364170 187398 364226
rect 187454 364170 187522 364226
rect 187578 364170 187648 364226
rect 187328 364102 187648 364170
rect 187328 364046 187398 364102
rect 187454 364046 187522 364102
rect 187578 364046 187648 364102
rect 187328 363978 187648 364046
rect 187328 363922 187398 363978
rect 187454 363922 187522 363978
rect 187578 363922 187648 363978
rect 187328 363888 187648 363922
rect 218048 364350 218368 364384
rect 218048 364294 218118 364350
rect 218174 364294 218242 364350
rect 218298 364294 218368 364350
rect 218048 364226 218368 364294
rect 218048 364170 218118 364226
rect 218174 364170 218242 364226
rect 218298 364170 218368 364226
rect 218048 364102 218368 364170
rect 218048 364046 218118 364102
rect 218174 364046 218242 364102
rect 218298 364046 218368 364102
rect 218048 363978 218368 364046
rect 218048 363922 218118 363978
rect 218174 363922 218242 363978
rect 218298 363922 218368 363978
rect 218048 363888 218368 363922
rect 248768 364350 249088 364384
rect 248768 364294 248838 364350
rect 248894 364294 248962 364350
rect 249018 364294 249088 364350
rect 248768 364226 249088 364294
rect 248768 364170 248838 364226
rect 248894 364170 248962 364226
rect 249018 364170 249088 364226
rect 248768 364102 249088 364170
rect 248768 364046 248838 364102
rect 248894 364046 248962 364102
rect 249018 364046 249088 364102
rect 248768 363978 249088 364046
rect 248768 363922 248838 363978
rect 248894 363922 248962 363978
rect 249018 363922 249088 363978
rect 248768 363888 249088 363922
rect 273084 363300 273140 363310
rect 110528 352350 110848 352384
rect 110528 352294 110598 352350
rect 110654 352294 110722 352350
rect 110778 352294 110848 352350
rect 110528 352226 110848 352294
rect 110528 352170 110598 352226
rect 110654 352170 110722 352226
rect 110778 352170 110848 352226
rect 110528 352102 110848 352170
rect 110528 352046 110598 352102
rect 110654 352046 110722 352102
rect 110778 352046 110848 352102
rect 110528 351978 110848 352046
rect 110528 351922 110598 351978
rect 110654 351922 110722 351978
rect 110778 351922 110848 351978
rect 110528 351888 110848 351922
rect 141248 352350 141568 352384
rect 141248 352294 141318 352350
rect 141374 352294 141442 352350
rect 141498 352294 141568 352350
rect 141248 352226 141568 352294
rect 141248 352170 141318 352226
rect 141374 352170 141442 352226
rect 141498 352170 141568 352226
rect 141248 352102 141568 352170
rect 141248 352046 141318 352102
rect 141374 352046 141442 352102
rect 141498 352046 141568 352102
rect 141248 351978 141568 352046
rect 141248 351922 141318 351978
rect 141374 351922 141442 351978
rect 141498 351922 141568 351978
rect 141248 351888 141568 351922
rect 171968 352350 172288 352384
rect 171968 352294 172038 352350
rect 172094 352294 172162 352350
rect 172218 352294 172288 352350
rect 171968 352226 172288 352294
rect 171968 352170 172038 352226
rect 172094 352170 172162 352226
rect 172218 352170 172288 352226
rect 171968 352102 172288 352170
rect 171968 352046 172038 352102
rect 172094 352046 172162 352102
rect 172218 352046 172288 352102
rect 171968 351978 172288 352046
rect 171968 351922 172038 351978
rect 172094 351922 172162 351978
rect 172218 351922 172288 351978
rect 171968 351888 172288 351922
rect 202688 352350 203008 352384
rect 202688 352294 202758 352350
rect 202814 352294 202882 352350
rect 202938 352294 203008 352350
rect 202688 352226 203008 352294
rect 202688 352170 202758 352226
rect 202814 352170 202882 352226
rect 202938 352170 203008 352226
rect 202688 352102 203008 352170
rect 202688 352046 202758 352102
rect 202814 352046 202882 352102
rect 202938 352046 203008 352102
rect 202688 351978 203008 352046
rect 202688 351922 202758 351978
rect 202814 351922 202882 351978
rect 202938 351922 203008 351978
rect 202688 351888 203008 351922
rect 233408 352350 233728 352384
rect 233408 352294 233478 352350
rect 233534 352294 233602 352350
rect 233658 352294 233728 352350
rect 233408 352226 233728 352294
rect 233408 352170 233478 352226
rect 233534 352170 233602 352226
rect 233658 352170 233728 352226
rect 233408 352102 233728 352170
rect 233408 352046 233478 352102
rect 233534 352046 233602 352102
rect 233658 352046 233728 352102
rect 233408 351978 233728 352046
rect 233408 351922 233478 351978
rect 233534 351922 233602 351978
rect 233658 351922 233728 351978
rect 233408 351888 233728 351922
rect 264128 352350 264448 352384
rect 264128 352294 264198 352350
rect 264254 352294 264322 352350
rect 264378 352294 264448 352350
rect 264128 352226 264448 352294
rect 264128 352170 264198 352226
rect 264254 352170 264322 352226
rect 264378 352170 264448 352226
rect 264128 352102 264448 352170
rect 264128 352046 264198 352102
rect 264254 352046 264322 352102
rect 264378 352046 264448 352102
rect 264128 351978 264448 352046
rect 264128 351922 264198 351978
rect 264254 351922 264322 351978
rect 264378 351922 264448 351978
rect 264128 351888 264448 351922
rect 95168 346350 95488 346384
rect 95168 346294 95238 346350
rect 95294 346294 95362 346350
rect 95418 346294 95488 346350
rect 95168 346226 95488 346294
rect 95168 346170 95238 346226
rect 95294 346170 95362 346226
rect 95418 346170 95488 346226
rect 95168 346102 95488 346170
rect 95168 346046 95238 346102
rect 95294 346046 95362 346102
rect 95418 346046 95488 346102
rect 95168 345978 95488 346046
rect 95168 345922 95238 345978
rect 95294 345922 95362 345978
rect 95418 345922 95488 345978
rect 95168 345888 95488 345922
rect 125888 346350 126208 346384
rect 125888 346294 125958 346350
rect 126014 346294 126082 346350
rect 126138 346294 126208 346350
rect 125888 346226 126208 346294
rect 125888 346170 125958 346226
rect 126014 346170 126082 346226
rect 126138 346170 126208 346226
rect 125888 346102 126208 346170
rect 125888 346046 125958 346102
rect 126014 346046 126082 346102
rect 126138 346046 126208 346102
rect 125888 345978 126208 346046
rect 125888 345922 125958 345978
rect 126014 345922 126082 345978
rect 126138 345922 126208 345978
rect 125888 345888 126208 345922
rect 156608 346350 156928 346384
rect 156608 346294 156678 346350
rect 156734 346294 156802 346350
rect 156858 346294 156928 346350
rect 156608 346226 156928 346294
rect 156608 346170 156678 346226
rect 156734 346170 156802 346226
rect 156858 346170 156928 346226
rect 156608 346102 156928 346170
rect 156608 346046 156678 346102
rect 156734 346046 156802 346102
rect 156858 346046 156928 346102
rect 156608 345978 156928 346046
rect 156608 345922 156678 345978
rect 156734 345922 156802 345978
rect 156858 345922 156928 345978
rect 156608 345888 156928 345922
rect 187328 346350 187648 346384
rect 187328 346294 187398 346350
rect 187454 346294 187522 346350
rect 187578 346294 187648 346350
rect 187328 346226 187648 346294
rect 187328 346170 187398 346226
rect 187454 346170 187522 346226
rect 187578 346170 187648 346226
rect 187328 346102 187648 346170
rect 187328 346046 187398 346102
rect 187454 346046 187522 346102
rect 187578 346046 187648 346102
rect 187328 345978 187648 346046
rect 187328 345922 187398 345978
rect 187454 345922 187522 345978
rect 187578 345922 187648 345978
rect 187328 345888 187648 345922
rect 218048 346350 218368 346384
rect 218048 346294 218118 346350
rect 218174 346294 218242 346350
rect 218298 346294 218368 346350
rect 218048 346226 218368 346294
rect 218048 346170 218118 346226
rect 218174 346170 218242 346226
rect 218298 346170 218368 346226
rect 218048 346102 218368 346170
rect 218048 346046 218118 346102
rect 218174 346046 218242 346102
rect 218298 346046 218368 346102
rect 218048 345978 218368 346046
rect 218048 345922 218118 345978
rect 218174 345922 218242 345978
rect 218298 345922 218368 345978
rect 218048 345888 218368 345922
rect 248768 346350 249088 346384
rect 248768 346294 248838 346350
rect 248894 346294 248962 346350
rect 249018 346294 249088 346350
rect 248768 346226 249088 346294
rect 248768 346170 248838 346226
rect 248894 346170 248962 346226
rect 249018 346170 249088 346226
rect 248768 346102 249088 346170
rect 248768 346046 248838 346102
rect 248894 346046 248962 346102
rect 249018 346046 249088 346102
rect 248768 345978 249088 346046
rect 248768 345922 248838 345978
rect 248894 345922 248962 345978
rect 249018 345922 249088 345978
rect 248768 345888 249088 345922
rect 272972 344484 273028 344494
rect 110528 334350 110848 334384
rect 110528 334294 110598 334350
rect 110654 334294 110722 334350
rect 110778 334294 110848 334350
rect 110528 334226 110848 334294
rect 110528 334170 110598 334226
rect 110654 334170 110722 334226
rect 110778 334170 110848 334226
rect 110528 334102 110848 334170
rect 110528 334046 110598 334102
rect 110654 334046 110722 334102
rect 110778 334046 110848 334102
rect 110528 333978 110848 334046
rect 110528 333922 110598 333978
rect 110654 333922 110722 333978
rect 110778 333922 110848 333978
rect 110528 333888 110848 333922
rect 141248 334350 141568 334384
rect 141248 334294 141318 334350
rect 141374 334294 141442 334350
rect 141498 334294 141568 334350
rect 141248 334226 141568 334294
rect 141248 334170 141318 334226
rect 141374 334170 141442 334226
rect 141498 334170 141568 334226
rect 141248 334102 141568 334170
rect 141248 334046 141318 334102
rect 141374 334046 141442 334102
rect 141498 334046 141568 334102
rect 141248 333978 141568 334046
rect 141248 333922 141318 333978
rect 141374 333922 141442 333978
rect 141498 333922 141568 333978
rect 141248 333888 141568 333922
rect 171968 334350 172288 334384
rect 171968 334294 172038 334350
rect 172094 334294 172162 334350
rect 172218 334294 172288 334350
rect 171968 334226 172288 334294
rect 171968 334170 172038 334226
rect 172094 334170 172162 334226
rect 172218 334170 172288 334226
rect 171968 334102 172288 334170
rect 171968 334046 172038 334102
rect 172094 334046 172162 334102
rect 172218 334046 172288 334102
rect 171968 333978 172288 334046
rect 171968 333922 172038 333978
rect 172094 333922 172162 333978
rect 172218 333922 172288 333978
rect 171968 333888 172288 333922
rect 202688 334350 203008 334384
rect 202688 334294 202758 334350
rect 202814 334294 202882 334350
rect 202938 334294 203008 334350
rect 202688 334226 203008 334294
rect 202688 334170 202758 334226
rect 202814 334170 202882 334226
rect 202938 334170 203008 334226
rect 202688 334102 203008 334170
rect 202688 334046 202758 334102
rect 202814 334046 202882 334102
rect 202938 334046 203008 334102
rect 202688 333978 203008 334046
rect 202688 333922 202758 333978
rect 202814 333922 202882 333978
rect 202938 333922 203008 333978
rect 202688 333888 203008 333922
rect 233408 334350 233728 334384
rect 233408 334294 233478 334350
rect 233534 334294 233602 334350
rect 233658 334294 233728 334350
rect 233408 334226 233728 334294
rect 233408 334170 233478 334226
rect 233534 334170 233602 334226
rect 233658 334170 233728 334226
rect 233408 334102 233728 334170
rect 233408 334046 233478 334102
rect 233534 334046 233602 334102
rect 233658 334046 233728 334102
rect 233408 333978 233728 334046
rect 233408 333922 233478 333978
rect 233534 333922 233602 333978
rect 233658 333922 233728 333978
rect 233408 333888 233728 333922
rect 264128 334350 264448 334384
rect 264128 334294 264198 334350
rect 264254 334294 264322 334350
rect 264378 334294 264448 334350
rect 264128 334226 264448 334294
rect 264128 334170 264198 334226
rect 264254 334170 264322 334226
rect 264378 334170 264448 334226
rect 264128 334102 264448 334170
rect 264128 334046 264198 334102
rect 264254 334046 264322 334102
rect 264378 334046 264448 334102
rect 264128 333978 264448 334046
rect 264128 333922 264198 333978
rect 264254 333922 264322 333978
rect 264378 333922 264448 333978
rect 264128 333888 264448 333922
rect 84812 300112 84868 300122
rect 84924 329338 84980 329348
rect 83804 298852 83860 298862
rect 84924 297298 84980 329282
rect 95168 328350 95488 328384
rect 95168 328294 95238 328350
rect 95294 328294 95362 328350
rect 95418 328294 95488 328350
rect 95168 328226 95488 328294
rect 95168 328170 95238 328226
rect 95294 328170 95362 328226
rect 95418 328170 95488 328226
rect 95168 328102 95488 328170
rect 95168 328046 95238 328102
rect 95294 328046 95362 328102
rect 95418 328046 95488 328102
rect 95168 327978 95488 328046
rect 95168 327922 95238 327978
rect 95294 327922 95362 327978
rect 95418 327922 95488 327978
rect 95168 327888 95488 327922
rect 125888 328350 126208 328384
rect 125888 328294 125958 328350
rect 126014 328294 126082 328350
rect 126138 328294 126208 328350
rect 125888 328226 126208 328294
rect 125888 328170 125958 328226
rect 126014 328170 126082 328226
rect 126138 328170 126208 328226
rect 125888 328102 126208 328170
rect 125888 328046 125958 328102
rect 126014 328046 126082 328102
rect 126138 328046 126208 328102
rect 125888 327978 126208 328046
rect 125888 327922 125958 327978
rect 126014 327922 126082 327978
rect 126138 327922 126208 327978
rect 125888 327888 126208 327922
rect 156608 328350 156928 328384
rect 156608 328294 156678 328350
rect 156734 328294 156802 328350
rect 156858 328294 156928 328350
rect 156608 328226 156928 328294
rect 156608 328170 156678 328226
rect 156734 328170 156802 328226
rect 156858 328170 156928 328226
rect 156608 328102 156928 328170
rect 156608 328046 156678 328102
rect 156734 328046 156802 328102
rect 156858 328046 156928 328102
rect 156608 327978 156928 328046
rect 156608 327922 156678 327978
rect 156734 327922 156802 327978
rect 156858 327922 156928 327978
rect 156608 327888 156928 327922
rect 187328 328350 187648 328384
rect 187328 328294 187398 328350
rect 187454 328294 187522 328350
rect 187578 328294 187648 328350
rect 187328 328226 187648 328294
rect 187328 328170 187398 328226
rect 187454 328170 187522 328226
rect 187578 328170 187648 328226
rect 187328 328102 187648 328170
rect 187328 328046 187398 328102
rect 187454 328046 187522 328102
rect 187578 328046 187648 328102
rect 187328 327978 187648 328046
rect 187328 327922 187398 327978
rect 187454 327922 187522 327978
rect 187578 327922 187648 327978
rect 187328 327888 187648 327922
rect 218048 328350 218368 328384
rect 218048 328294 218118 328350
rect 218174 328294 218242 328350
rect 218298 328294 218368 328350
rect 218048 328226 218368 328294
rect 218048 328170 218118 328226
rect 218174 328170 218242 328226
rect 218298 328170 218368 328226
rect 218048 328102 218368 328170
rect 218048 328046 218118 328102
rect 218174 328046 218242 328102
rect 218298 328046 218368 328102
rect 218048 327978 218368 328046
rect 218048 327922 218118 327978
rect 218174 327922 218242 327978
rect 218298 327922 218368 327978
rect 218048 327888 218368 327922
rect 248768 328350 249088 328384
rect 248768 328294 248838 328350
rect 248894 328294 248962 328350
rect 249018 328294 249088 328350
rect 248768 328226 249088 328294
rect 248768 328170 248838 328226
rect 248894 328170 248962 328226
rect 249018 328170 249088 328226
rect 248768 328102 249088 328170
rect 248768 328046 248838 328102
rect 248894 328046 248962 328102
rect 249018 328046 249088 328102
rect 248768 327978 249088 328046
rect 248768 327922 248838 327978
rect 248894 327922 248962 327978
rect 249018 327922 249088 327978
rect 248768 327888 249088 327922
rect 272972 319978 273028 344428
rect 273084 343558 273140 363244
rect 273756 361956 273812 361966
rect 273756 361378 273812 361900
rect 273756 361312 273812 361322
rect 273756 360612 273812 360622
rect 273308 359268 273364 359278
rect 273308 350218 273364 359212
rect 273756 358678 273812 360556
rect 273756 358612 273812 358622
rect 273644 357924 273700 357934
rect 273644 353638 273700 357868
rect 273756 356580 273812 356590
rect 273756 356338 273812 356524
rect 273756 356272 273812 356282
rect 273756 355236 273812 355246
rect 273756 354538 273812 355180
rect 273756 354472 273812 354482
rect 273756 353638 273812 353648
rect 273644 353582 273756 353638
rect 273756 353572 273812 353582
rect 273308 350152 273364 350162
rect 273644 351204 273700 351214
rect 273084 343492 273140 343502
rect 273644 341938 273700 351148
rect 273756 349860 273812 349870
rect 273756 349498 273812 349804
rect 273756 349432 273812 349442
rect 273756 348516 273812 348526
rect 273756 343738 273812 348460
rect 273756 343672 273812 343682
rect 273644 341872 273700 341882
rect 273196 341796 273252 341806
rect 272972 319912 273028 319922
rect 273084 336420 273140 336430
rect 110528 316350 110848 316384
rect 110528 316294 110598 316350
rect 110654 316294 110722 316350
rect 110778 316294 110848 316350
rect 110528 316226 110848 316294
rect 110528 316170 110598 316226
rect 110654 316170 110722 316226
rect 110778 316170 110848 316226
rect 110528 316102 110848 316170
rect 110528 316046 110598 316102
rect 110654 316046 110722 316102
rect 110778 316046 110848 316102
rect 110528 315978 110848 316046
rect 110528 315922 110598 315978
rect 110654 315922 110722 315978
rect 110778 315922 110848 315978
rect 110528 315888 110848 315922
rect 141248 316350 141568 316384
rect 141248 316294 141318 316350
rect 141374 316294 141442 316350
rect 141498 316294 141568 316350
rect 141248 316226 141568 316294
rect 141248 316170 141318 316226
rect 141374 316170 141442 316226
rect 141498 316170 141568 316226
rect 141248 316102 141568 316170
rect 141248 316046 141318 316102
rect 141374 316046 141442 316102
rect 141498 316046 141568 316102
rect 141248 315978 141568 316046
rect 141248 315922 141318 315978
rect 141374 315922 141442 315978
rect 141498 315922 141568 315978
rect 141248 315888 141568 315922
rect 171968 316350 172288 316384
rect 171968 316294 172038 316350
rect 172094 316294 172162 316350
rect 172218 316294 172288 316350
rect 171968 316226 172288 316294
rect 171968 316170 172038 316226
rect 172094 316170 172162 316226
rect 172218 316170 172288 316226
rect 171968 316102 172288 316170
rect 171968 316046 172038 316102
rect 172094 316046 172162 316102
rect 172218 316046 172288 316102
rect 171968 315978 172288 316046
rect 171968 315922 172038 315978
rect 172094 315922 172162 315978
rect 172218 315922 172288 315978
rect 171968 315888 172288 315922
rect 202688 316350 203008 316384
rect 202688 316294 202758 316350
rect 202814 316294 202882 316350
rect 202938 316294 203008 316350
rect 202688 316226 203008 316294
rect 202688 316170 202758 316226
rect 202814 316170 202882 316226
rect 202938 316170 203008 316226
rect 202688 316102 203008 316170
rect 202688 316046 202758 316102
rect 202814 316046 202882 316102
rect 202938 316046 203008 316102
rect 202688 315978 203008 316046
rect 202688 315922 202758 315978
rect 202814 315922 202882 315978
rect 202938 315922 203008 315978
rect 202688 315888 203008 315922
rect 233408 316350 233728 316384
rect 233408 316294 233478 316350
rect 233534 316294 233602 316350
rect 233658 316294 233728 316350
rect 233408 316226 233728 316294
rect 233408 316170 233478 316226
rect 233534 316170 233602 316226
rect 233658 316170 233728 316226
rect 233408 316102 233728 316170
rect 233408 316046 233478 316102
rect 233534 316046 233602 316102
rect 233658 316046 233728 316102
rect 233408 315978 233728 316046
rect 233408 315922 233478 315978
rect 233534 315922 233602 315978
rect 233658 315922 233728 315978
rect 233408 315888 233728 315922
rect 264128 316350 264448 316384
rect 264128 316294 264198 316350
rect 264254 316294 264322 316350
rect 264378 316294 264448 316350
rect 264128 316226 264448 316294
rect 264128 316170 264198 316226
rect 264254 316170 264322 316226
rect 264378 316170 264448 316226
rect 264128 316102 264448 316170
rect 264128 316046 264198 316102
rect 264254 316046 264322 316102
rect 264378 316046 264448 316102
rect 264128 315978 264448 316046
rect 264128 315922 264198 315978
rect 264254 315922 264322 315978
rect 264378 315922 264448 315978
rect 264128 315888 264448 315922
rect 273084 311698 273140 336364
rect 273196 323398 273252 341740
rect 273756 340452 273812 340462
rect 273308 337764 273364 337774
rect 273308 325018 273364 337708
rect 273756 330058 273812 340396
rect 278012 333658 278068 430556
rect 278124 430052 278180 430062
rect 278124 335998 278180 429996
rect 279692 429156 279748 429166
rect 278124 335932 278180 335942
rect 278236 376498 278292 376508
rect 278012 333592 278068 333602
rect 273756 329992 273812 330002
rect 273308 324952 273364 324962
rect 273196 323332 273252 323342
rect 273084 311632 273140 311642
rect 274652 317638 274708 317648
rect 272188 310884 272244 310894
rect 95168 310350 95488 310384
rect 95168 310294 95238 310350
rect 95294 310294 95362 310350
rect 95418 310294 95488 310350
rect 95168 310226 95488 310294
rect 95168 310170 95238 310226
rect 95294 310170 95362 310226
rect 95418 310170 95488 310226
rect 95168 310102 95488 310170
rect 95168 310046 95238 310102
rect 95294 310046 95362 310102
rect 95418 310046 95488 310102
rect 95168 309978 95488 310046
rect 95168 309922 95238 309978
rect 95294 309922 95362 309978
rect 95418 309922 95488 309978
rect 95168 309888 95488 309922
rect 125888 310350 126208 310384
rect 125888 310294 125958 310350
rect 126014 310294 126082 310350
rect 126138 310294 126208 310350
rect 125888 310226 126208 310294
rect 125888 310170 125958 310226
rect 126014 310170 126082 310226
rect 126138 310170 126208 310226
rect 125888 310102 126208 310170
rect 125888 310046 125958 310102
rect 126014 310046 126082 310102
rect 126138 310046 126208 310102
rect 125888 309978 126208 310046
rect 125888 309922 125958 309978
rect 126014 309922 126082 309978
rect 126138 309922 126208 309978
rect 125888 309888 126208 309922
rect 156608 310350 156928 310384
rect 156608 310294 156678 310350
rect 156734 310294 156802 310350
rect 156858 310294 156928 310350
rect 156608 310226 156928 310294
rect 156608 310170 156678 310226
rect 156734 310170 156802 310226
rect 156858 310170 156928 310226
rect 156608 310102 156928 310170
rect 156608 310046 156678 310102
rect 156734 310046 156802 310102
rect 156858 310046 156928 310102
rect 156608 309978 156928 310046
rect 156608 309922 156678 309978
rect 156734 309922 156802 309978
rect 156858 309922 156928 309978
rect 156608 309888 156928 309922
rect 187328 310350 187648 310384
rect 187328 310294 187398 310350
rect 187454 310294 187522 310350
rect 187578 310294 187648 310350
rect 187328 310226 187648 310294
rect 187328 310170 187398 310226
rect 187454 310170 187522 310226
rect 187578 310170 187648 310226
rect 187328 310102 187648 310170
rect 187328 310046 187398 310102
rect 187454 310046 187522 310102
rect 187578 310046 187648 310102
rect 187328 309978 187648 310046
rect 187328 309922 187398 309978
rect 187454 309922 187522 309978
rect 187578 309922 187648 309978
rect 187328 309888 187648 309922
rect 218048 310350 218368 310384
rect 218048 310294 218118 310350
rect 218174 310294 218242 310350
rect 218298 310294 218368 310350
rect 218048 310226 218368 310294
rect 218048 310170 218118 310226
rect 218174 310170 218242 310226
rect 218298 310170 218368 310226
rect 218048 310102 218368 310170
rect 218048 310046 218118 310102
rect 218174 310046 218242 310102
rect 218298 310046 218368 310102
rect 218048 309978 218368 310046
rect 218048 309922 218118 309978
rect 218174 309922 218242 309978
rect 218298 309922 218368 309978
rect 218048 309888 218368 309922
rect 248768 310350 249088 310384
rect 248768 310294 248838 310350
rect 248894 310294 248962 310350
rect 249018 310294 249088 310350
rect 248768 310226 249088 310294
rect 248768 310170 248838 310226
rect 248894 310170 248962 310226
rect 249018 310170 249088 310226
rect 248768 310102 249088 310170
rect 248768 310046 248838 310102
rect 248894 310046 248962 310102
rect 249018 310046 249088 310102
rect 248768 309978 249088 310046
rect 248768 309922 248838 309978
rect 248894 309922 248962 309978
rect 249018 309922 249088 309978
rect 248768 309888 249088 309922
rect 84924 297232 84980 297242
rect 83692 295072 83748 295082
rect 83356 280354 83412 280364
rect 97578 292350 98198 299890
rect 97578 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 98198 292350
rect 97578 292226 98198 292294
rect 97578 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 98198 292226
rect 97578 292102 98198 292170
rect 97578 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 98198 292102
rect 97578 291978 98198 292046
rect 97578 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 98198 291978
rect 97578 274350 98198 291922
rect 97578 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 98198 274350
rect 97578 274226 98198 274294
rect 97578 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 98198 274226
rect 97578 274102 98198 274170
rect 97578 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 98198 274102
rect 97578 273978 98198 274046
rect 97578 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 98198 273978
rect 86492 258020 86548 258030
rect 84924 142324 84980 142334
rect 84924 142138 84980 142268
rect 84924 142072 84980 142082
rect 81452 4274 81508 4284
rect 80556 4162 80612 4172
rect 86492 4228 86548 257964
rect 97578 256350 98198 273922
rect 97578 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 98198 256350
rect 97578 256226 98198 256294
rect 97578 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 98198 256226
rect 97578 256102 98198 256170
rect 97578 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 98198 256102
rect 97578 255978 98198 256046
rect 97578 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 98198 255978
rect 97578 238350 98198 255922
rect 97578 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 98198 238350
rect 97578 238226 98198 238294
rect 97578 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 98198 238226
rect 97578 238102 98198 238170
rect 97578 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 98198 238102
rect 97578 237978 98198 238046
rect 97578 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 98198 237978
rect 89852 231140 89908 231150
rect 89852 4340 89908 231084
rect 97578 220350 98198 237922
rect 97578 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 98198 220350
rect 97578 220226 98198 220294
rect 97578 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 98198 220226
rect 97578 220102 98198 220170
rect 97578 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 98198 220102
rect 97578 219978 98198 220046
rect 97578 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 98198 219978
rect 95168 202350 95488 202384
rect 95168 202294 95238 202350
rect 95294 202294 95362 202350
rect 95418 202294 95488 202350
rect 95168 202226 95488 202294
rect 95168 202170 95238 202226
rect 95294 202170 95362 202226
rect 95418 202170 95488 202226
rect 95168 202102 95488 202170
rect 95168 202046 95238 202102
rect 95294 202046 95362 202102
rect 95418 202046 95488 202102
rect 95168 201978 95488 202046
rect 95168 201922 95238 201978
rect 95294 201922 95362 201978
rect 95418 201922 95488 201978
rect 95168 201888 95488 201922
rect 97578 202350 98198 219922
rect 97578 202294 97674 202350
rect 97730 202294 97798 202350
rect 97854 202294 97922 202350
rect 97978 202294 98046 202350
rect 98102 202294 98198 202350
rect 97578 202226 98198 202294
rect 97578 202170 97674 202226
rect 97730 202170 97798 202226
rect 97854 202170 97922 202226
rect 97978 202170 98046 202226
rect 98102 202170 98198 202226
rect 97578 202102 98198 202170
rect 97578 202046 97674 202102
rect 97730 202046 97798 202102
rect 97854 202046 97922 202102
rect 97978 202046 98046 202102
rect 98102 202046 98198 202102
rect 97578 201978 98198 202046
rect 97578 201922 97674 201978
rect 97730 201922 97798 201978
rect 97854 201922 97922 201978
rect 97978 201922 98046 201978
rect 98102 201922 98198 201978
rect 95168 184350 95488 184384
rect 95168 184294 95238 184350
rect 95294 184294 95362 184350
rect 95418 184294 95488 184350
rect 95168 184226 95488 184294
rect 95168 184170 95238 184226
rect 95294 184170 95362 184226
rect 95418 184170 95488 184226
rect 95168 184102 95488 184170
rect 95168 184046 95238 184102
rect 95294 184046 95362 184102
rect 95418 184046 95488 184102
rect 95168 183978 95488 184046
rect 95168 183922 95238 183978
rect 95294 183922 95362 183978
rect 95418 183922 95488 183978
rect 95168 183888 95488 183922
rect 97578 184350 98198 201922
rect 97578 184294 97674 184350
rect 97730 184294 97798 184350
rect 97854 184294 97922 184350
rect 97978 184294 98046 184350
rect 98102 184294 98198 184350
rect 97578 184226 98198 184294
rect 97578 184170 97674 184226
rect 97730 184170 97798 184226
rect 97854 184170 97922 184226
rect 97978 184170 98046 184226
rect 98102 184170 98198 184226
rect 97578 184102 98198 184170
rect 97578 184046 97674 184102
rect 97730 184046 97798 184102
rect 97854 184046 97922 184102
rect 97978 184046 98046 184102
rect 98102 184046 98198 184102
rect 97578 183978 98198 184046
rect 97578 183922 97674 183978
rect 97730 183922 97798 183978
rect 97854 183922 97922 183978
rect 97978 183922 98046 183978
rect 98102 183922 98198 183978
rect 95168 166350 95488 166384
rect 95168 166294 95238 166350
rect 95294 166294 95362 166350
rect 95418 166294 95488 166350
rect 95168 166226 95488 166294
rect 95168 166170 95238 166226
rect 95294 166170 95362 166226
rect 95418 166170 95488 166226
rect 95168 166102 95488 166170
rect 95168 166046 95238 166102
rect 95294 166046 95362 166102
rect 95418 166046 95488 166102
rect 95168 165978 95488 166046
rect 95168 165922 95238 165978
rect 95294 165922 95362 165978
rect 95418 165922 95488 165978
rect 95168 165888 95488 165922
rect 97578 166350 98198 183922
rect 97578 166294 97674 166350
rect 97730 166294 97798 166350
rect 97854 166294 97922 166350
rect 97978 166294 98046 166350
rect 98102 166294 98198 166350
rect 97578 166226 98198 166294
rect 97578 166170 97674 166226
rect 97730 166170 97798 166226
rect 97854 166170 97922 166226
rect 97978 166170 98046 166226
rect 98102 166170 98198 166226
rect 97578 166102 98198 166170
rect 97578 166046 97674 166102
rect 97730 166046 97798 166102
rect 97854 166046 97922 166102
rect 97978 166046 98046 166102
rect 98102 166046 98198 166102
rect 97578 165978 98198 166046
rect 97578 165922 97674 165978
rect 97730 165922 97798 165978
rect 97854 165922 97922 165978
rect 97978 165922 98046 165978
rect 98102 165922 98198 165978
rect 89852 4274 89908 4284
rect 97578 148350 98198 165922
rect 97578 148294 97674 148350
rect 97730 148294 97798 148350
rect 97854 148294 97922 148350
rect 97978 148294 98046 148350
rect 98102 148294 98198 148350
rect 97578 148226 98198 148294
rect 97578 148170 97674 148226
rect 97730 148170 97798 148226
rect 97854 148170 97922 148226
rect 97978 148170 98046 148226
rect 98102 148170 98198 148226
rect 97578 148102 98198 148170
rect 97578 148046 97674 148102
rect 97730 148046 97798 148102
rect 97854 148046 97922 148102
rect 97978 148046 98046 148102
rect 98102 148046 98198 148102
rect 97578 147978 98198 148046
rect 97578 147922 97674 147978
rect 97730 147922 97798 147978
rect 97854 147922 97922 147978
rect 97978 147922 98046 147978
rect 98102 147922 98198 147978
rect 97578 130350 98198 147922
rect 97578 130294 97674 130350
rect 97730 130294 97798 130350
rect 97854 130294 97922 130350
rect 97978 130294 98046 130350
rect 98102 130294 98198 130350
rect 97578 130226 98198 130294
rect 97578 130170 97674 130226
rect 97730 130170 97798 130226
rect 97854 130170 97922 130226
rect 97978 130170 98046 130226
rect 98102 130170 98198 130226
rect 97578 130102 98198 130170
rect 97578 130046 97674 130102
rect 97730 130046 97798 130102
rect 97854 130046 97922 130102
rect 97978 130046 98046 130102
rect 98102 130046 98198 130102
rect 97578 129978 98198 130046
rect 97578 129922 97674 129978
rect 97730 129922 97798 129978
rect 97854 129922 97922 129978
rect 97978 129922 98046 129978
rect 98102 129922 98198 129978
rect 97578 112350 98198 129922
rect 97578 112294 97674 112350
rect 97730 112294 97798 112350
rect 97854 112294 97922 112350
rect 97978 112294 98046 112350
rect 98102 112294 98198 112350
rect 97578 112226 98198 112294
rect 97578 112170 97674 112226
rect 97730 112170 97798 112226
rect 97854 112170 97922 112226
rect 97978 112170 98046 112226
rect 98102 112170 98198 112226
rect 97578 112102 98198 112170
rect 97578 112046 97674 112102
rect 97730 112046 97798 112102
rect 97854 112046 97922 112102
rect 97978 112046 98046 112102
rect 98102 112046 98198 112102
rect 97578 111978 98198 112046
rect 97578 111922 97674 111978
rect 97730 111922 97798 111978
rect 97854 111922 97922 111978
rect 97978 111922 98046 111978
rect 98102 111922 98198 111978
rect 97578 94350 98198 111922
rect 97578 94294 97674 94350
rect 97730 94294 97798 94350
rect 97854 94294 97922 94350
rect 97978 94294 98046 94350
rect 98102 94294 98198 94350
rect 97578 94226 98198 94294
rect 97578 94170 97674 94226
rect 97730 94170 97798 94226
rect 97854 94170 97922 94226
rect 97978 94170 98046 94226
rect 98102 94170 98198 94226
rect 97578 94102 98198 94170
rect 97578 94046 97674 94102
rect 97730 94046 97798 94102
rect 97854 94046 97922 94102
rect 97978 94046 98046 94102
rect 98102 94046 98198 94102
rect 97578 93978 98198 94046
rect 97578 93922 97674 93978
rect 97730 93922 97798 93978
rect 97854 93922 97922 93978
rect 97978 93922 98046 93978
rect 98102 93922 98198 93978
rect 97578 76350 98198 93922
rect 97578 76294 97674 76350
rect 97730 76294 97798 76350
rect 97854 76294 97922 76350
rect 97978 76294 98046 76350
rect 98102 76294 98198 76350
rect 97578 76226 98198 76294
rect 97578 76170 97674 76226
rect 97730 76170 97798 76226
rect 97854 76170 97922 76226
rect 97978 76170 98046 76226
rect 98102 76170 98198 76226
rect 97578 76102 98198 76170
rect 97578 76046 97674 76102
rect 97730 76046 97798 76102
rect 97854 76046 97922 76102
rect 97978 76046 98046 76102
rect 98102 76046 98198 76102
rect 97578 75978 98198 76046
rect 97578 75922 97674 75978
rect 97730 75922 97798 75978
rect 97854 75922 97922 75978
rect 97978 75922 98046 75978
rect 98102 75922 98198 75978
rect 97578 58350 98198 75922
rect 97578 58294 97674 58350
rect 97730 58294 97798 58350
rect 97854 58294 97922 58350
rect 97978 58294 98046 58350
rect 98102 58294 98198 58350
rect 97578 58226 98198 58294
rect 97578 58170 97674 58226
rect 97730 58170 97798 58226
rect 97854 58170 97922 58226
rect 97978 58170 98046 58226
rect 98102 58170 98198 58226
rect 97578 58102 98198 58170
rect 97578 58046 97674 58102
rect 97730 58046 97798 58102
rect 97854 58046 97922 58102
rect 97978 58046 98046 58102
rect 98102 58046 98198 58102
rect 97578 57978 98198 58046
rect 97578 57922 97674 57978
rect 97730 57922 97798 57978
rect 97854 57922 97922 57978
rect 97978 57922 98046 57978
rect 98102 57922 98198 57978
rect 97578 40350 98198 57922
rect 97578 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 98198 40350
rect 97578 40226 98198 40294
rect 97578 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 98198 40226
rect 97578 40102 98198 40170
rect 97578 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 98198 40102
rect 97578 39978 98198 40046
rect 97578 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 98198 39978
rect 97578 22350 98198 39922
rect 97578 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 98198 22350
rect 97578 22226 98198 22294
rect 97578 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 98198 22226
rect 97578 22102 98198 22170
rect 97578 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 98198 22102
rect 97578 21978 98198 22046
rect 97578 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 98198 21978
rect 97578 4350 98198 21922
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 86492 4162 86548 4172
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 298350 101918 299890
rect 101298 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 101918 298350
rect 101298 298226 101918 298294
rect 101298 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 101918 298226
rect 101298 298102 101918 298170
rect 101298 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 101918 298102
rect 101298 297978 101918 298046
rect 101298 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 101918 297978
rect 101298 280350 101918 297922
rect 110528 298350 110848 298384
rect 110528 298294 110598 298350
rect 110654 298294 110722 298350
rect 110778 298294 110848 298350
rect 110528 298226 110848 298294
rect 110528 298170 110598 298226
rect 110654 298170 110722 298226
rect 110778 298170 110848 298226
rect 110528 298102 110848 298170
rect 110528 298046 110598 298102
rect 110654 298046 110722 298102
rect 110778 298046 110848 298102
rect 110528 297978 110848 298046
rect 110528 297922 110598 297978
rect 110654 297922 110722 297978
rect 110778 297922 110848 297978
rect 110528 297888 110848 297922
rect 128298 292350 128918 299890
rect 128298 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 128918 292350
rect 128298 292226 128918 292294
rect 128298 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 128918 292226
rect 128298 292102 128918 292170
rect 128298 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 128918 292102
rect 128298 291978 128918 292046
rect 128298 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 128918 291978
rect 121772 286580 121828 286590
rect 101298 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 101918 280350
rect 101298 280226 101918 280294
rect 101298 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 101918 280226
rect 101298 280102 101918 280170
rect 101298 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 101918 280102
rect 101298 279978 101918 280046
rect 101298 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 101918 279978
rect 101298 262350 101918 279922
rect 101298 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 101918 262350
rect 101298 262226 101918 262294
rect 101298 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 101918 262226
rect 101298 262102 101918 262170
rect 101298 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 101918 262102
rect 101298 261978 101918 262046
rect 101298 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 101918 261978
rect 101298 244350 101918 261922
rect 101298 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 101918 244350
rect 101298 244226 101918 244294
rect 101298 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 101918 244226
rect 101298 244102 101918 244170
rect 101298 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 101918 244102
rect 101298 243978 101918 244046
rect 101298 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 101918 243978
rect 101298 226350 101918 243922
rect 101298 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 101918 226350
rect 101298 226226 101918 226294
rect 101298 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 101918 226226
rect 101298 226102 101918 226170
rect 101298 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 101918 226102
rect 101298 225978 101918 226046
rect 101298 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 101918 225978
rect 101298 208350 101918 225922
rect 101298 208294 101394 208350
rect 101450 208294 101518 208350
rect 101574 208294 101642 208350
rect 101698 208294 101766 208350
rect 101822 208294 101918 208350
rect 101298 208226 101918 208294
rect 101298 208170 101394 208226
rect 101450 208170 101518 208226
rect 101574 208170 101642 208226
rect 101698 208170 101766 208226
rect 101822 208170 101918 208226
rect 101298 208102 101918 208170
rect 101298 208046 101394 208102
rect 101450 208046 101518 208102
rect 101574 208046 101642 208102
rect 101698 208046 101766 208102
rect 101822 208046 101918 208102
rect 101298 207978 101918 208046
rect 101298 207922 101394 207978
rect 101450 207922 101518 207978
rect 101574 207922 101642 207978
rect 101698 207922 101766 207978
rect 101822 207922 101918 207978
rect 101298 190350 101918 207922
rect 101298 190294 101394 190350
rect 101450 190294 101518 190350
rect 101574 190294 101642 190350
rect 101698 190294 101766 190350
rect 101822 190294 101918 190350
rect 101298 190226 101918 190294
rect 101298 190170 101394 190226
rect 101450 190170 101518 190226
rect 101574 190170 101642 190226
rect 101698 190170 101766 190226
rect 101822 190170 101918 190226
rect 101298 190102 101918 190170
rect 101298 190046 101394 190102
rect 101450 190046 101518 190102
rect 101574 190046 101642 190102
rect 101698 190046 101766 190102
rect 101822 190046 101918 190102
rect 101298 189978 101918 190046
rect 101298 189922 101394 189978
rect 101450 189922 101518 189978
rect 101574 189922 101642 189978
rect 101698 189922 101766 189978
rect 101822 189922 101918 189978
rect 101298 172350 101918 189922
rect 101298 172294 101394 172350
rect 101450 172294 101518 172350
rect 101574 172294 101642 172350
rect 101698 172294 101766 172350
rect 101822 172294 101918 172350
rect 101298 172226 101918 172294
rect 101298 172170 101394 172226
rect 101450 172170 101518 172226
rect 101574 172170 101642 172226
rect 101698 172170 101766 172226
rect 101822 172170 101918 172226
rect 101298 172102 101918 172170
rect 101298 172046 101394 172102
rect 101450 172046 101518 172102
rect 101574 172046 101642 172102
rect 101698 172046 101766 172102
rect 101822 172046 101918 172102
rect 101298 171978 101918 172046
rect 101298 171922 101394 171978
rect 101450 171922 101518 171978
rect 101574 171922 101642 171978
rect 101698 171922 101766 171978
rect 101822 171922 101918 171978
rect 101298 154350 101918 171922
rect 101298 154294 101394 154350
rect 101450 154294 101518 154350
rect 101574 154294 101642 154350
rect 101698 154294 101766 154350
rect 101822 154294 101918 154350
rect 101298 154226 101918 154294
rect 101298 154170 101394 154226
rect 101450 154170 101518 154226
rect 101574 154170 101642 154226
rect 101698 154170 101766 154226
rect 101822 154170 101918 154226
rect 101298 154102 101918 154170
rect 101298 154046 101394 154102
rect 101450 154046 101518 154102
rect 101574 154046 101642 154102
rect 101698 154046 101766 154102
rect 101822 154046 101918 154102
rect 101298 153978 101918 154046
rect 101298 153922 101394 153978
rect 101450 153922 101518 153978
rect 101574 153922 101642 153978
rect 101698 153922 101766 153978
rect 101822 153922 101918 153978
rect 101298 136350 101918 153922
rect 101298 136294 101394 136350
rect 101450 136294 101518 136350
rect 101574 136294 101642 136350
rect 101698 136294 101766 136350
rect 101822 136294 101918 136350
rect 101298 136226 101918 136294
rect 101298 136170 101394 136226
rect 101450 136170 101518 136226
rect 101574 136170 101642 136226
rect 101698 136170 101766 136226
rect 101822 136170 101918 136226
rect 101298 136102 101918 136170
rect 101298 136046 101394 136102
rect 101450 136046 101518 136102
rect 101574 136046 101642 136102
rect 101698 136046 101766 136102
rect 101822 136046 101918 136102
rect 101298 135978 101918 136046
rect 101298 135922 101394 135978
rect 101450 135922 101518 135978
rect 101574 135922 101642 135978
rect 101698 135922 101766 135978
rect 101822 135922 101918 135978
rect 101298 118350 101918 135922
rect 101298 118294 101394 118350
rect 101450 118294 101518 118350
rect 101574 118294 101642 118350
rect 101698 118294 101766 118350
rect 101822 118294 101918 118350
rect 101298 118226 101918 118294
rect 101298 118170 101394 118226
rect 101450 118170 101518 118226
rect 101574 118170 101642 118226
rect 101698 118170 101766 118226
rect 101822 118170 101918 118226
rect 101298 118102 101918 118170
rect 101298 118046 101394 118102
rect 101450 118046 101518 118102
rect 101574 118046 101642 118102
rect 101698 118046 101766 118102
rect 101822 118046 101918 118102
rect 101298 117978 101918 118046
rect 101298 117922 101394 117978
rect 101450 117922 101518 117978
rect 101574 117922 101642 117978
rect 101698 117922 101766 117978
rect 101822 117922 101918 117978
rect 101298 100350 101918 117922
rect 101298 100294 101394 100350
rect 101450 100294 101518 100350
rect 101574 100294 101642 100350
rect 101698 100294 101766 100350
rect 101822 100294 101918 100350
rect 101298 100226 101918 100294
rect 101298 100170 101394 100226
rect 101450 100170 101518 100226
rect 101574 100170 101642 100226
rect 101698 100170 101766 100226
rect 101822 100170 101918 100226
rect 101298 100102 101918 100170
rect 101298 100046 101394 100102
rect 101450 100046 101518 100102
rect 101574 100046 101642 100102
rect 101698 100046 101766 100102
rect 101822 100046 101918 100102
rect 101298 99978 101918 100046
rect 101298 99922 101394 99978
rect 101450 99922 101518 99978
rect 101574 99922 101642 99978
rect 101698 99922 101766 99978
rect 101822 99922 101918 99978
rect 101298 82350 101918 99922
rect 101298 82294 101394 82350
rect 101450 82294 101518 82350
rect 101574 82294 101642 82350
rect 101698 82294 101766 82350
rect 101822 82294 101918 82350
rect 101298 82226 101918 82294
rect 101298 82170 101394 82226
rect 101450 82170 101518 82226
rect 101574 82170 101642 82226
rect 101698 82170 101766 82226
rect 101822 82170 101918 82226
rect 101298 82102 101918 82170
rect 101298 82046 101394 82102
rect 101450 82046 101518 82102
rect 101574 82046 101642 82102
rect 101698 82046 101766 82102
rect 101822 82046 101918 82102
rect 101298 81978 101918 82046
rect 101298 81922 101394 81978
rect 101450 81922 101518 81978
rect 101574 81922 101642 81978
rect 101698 81922 101766 81978
rect 101822 81922 101918 81978
rect 101298 64350 101918 81922
rect 101298 64294 101394 64350
rect 101450 64294 101518 64350
rect 101574 64294 101642 64350
rect 101698 64294 101766 64350
rect 101822 64294 101918 64350
rect 101298 64226 101918 64294
rect 101298 64170 101394 64226
rect 101450 64170 101518 64226
rect 101574 64170 101642 64226
rect 101698 64170 101766 64226
rect 101822 64170 101918 64226
rect 101298 64102 101918 64170
rect 101298 64046 101394 64102
rect 101450 64046 101518 64102
rect 101574 64046 101642 64102
rect 101698 64046 101766 64102
rect 101822 64046 101918 64102
rect 101298 63978 101918 64046
rect 101298 63922 101394 63978
rect 101450 63922 101518 63978
rect 101574 63922 101642 63978
rect 101698 63922 101766 63978
rect 101822 63922 101918 63978
rect 101298 46350 101918 63922
rect 101298 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 101918 46350
rect 101298 46226 101918 46294
rect 101298 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 101918 46226
rect 101298 46102 101918 46170
rect 101298 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 101918 46102
rect 101298 45978 101918 46046
rect 101298 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 101918 45978
rect 101298 28350 101918 45922
rect 101298 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 101918 28350
rect 101298 28226 101918 28294
rect 101298 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 101918 28226
rect 101298 28102 101918 28170
rect 101298 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 101918 28102
rect 101298 27978 101918 28046
rect 101298 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 101918 27978
rect 101298 10350 101918 27922
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 101298 -1120 101918 9922
rect 104972 285124 105028 285134
rect 104972 4228 105028 285068
rect 116732 283332 116788 283342
rect 104972 4162 105028 4172
rect 109116 222628 109172 222638
rect 109116 4228 109172 222572
rect 112476 209412 112532 209422
rect 110528 190350 110848 190384
rect 110528 190294 110598 190350
rect 110654 190294 110722 190350
rect 110778 190294 110848 190350
rect 110528 190226 110848 190294
rect 110528 190170 110598 190226
rect 110654 190170 110722 190226
rect 110778 190170 110848 190226
rect 110528 190102 110848 190170
rect 110528 190046 110598 190102
rect 110654 190046 110722 190102
rect 110778 190046 110848 190102
rect 110528 189978 110848 190046
rect 110528 189922 110598 189978
rect 110654 189922 110722 189978
rect 110778 189922 110848 189978
rect 110528 189888 110848 189922
rect 110528 172350 110848 172384
rect 110528 172294 110598 172350
rect 110654 172294 110722 172350
rect 110778 172294 110848 172350
rect 110528 172226 110848 172294
rect 110528 172170 110598 172226
rect 110654 172170 110722 172226
rect 110778 172170 110848 172226
rect 110528 172102 110848 172170
rect 110528 172046 110598 172102
rect 110654 172046 110722 172102
rect 110778 172046 110848 172102
rect 110528 171978 110848 172046
rect 110528 171922 110598 171978
rect 110654 171922 110722 171978
rect 110778 171922 110848 171978
rect 110528 171888 110848 171922
rect 109116 4162 109172 4172
rect 112476 4228 112532 209356
rect 114716 145572 114772 145582
rect 114716 141204 114772 145516
rect 114716 141058 114772 141148
rect 114716 140992 114772 141002
rect 112476 4162 112532 4172
rect 116732 4228 116788 283276
rect 116732 4162 116788 4172
rect 119196 210868 119252 210878
rect 119196 4228 119252 210812
rect 119308 142678 119364 142688
rect 119308 141958 119364 142622
rect 119308 141204 119364 141902
rect 119308 141138 119364 141148
rect 121772 26068 121828 286524
rect 123452 286356 123508 286366
rect 123452 158900 123508 286300
rect 123452 158834 123508 158844
rect 124348 285684 124404 285694
rect 124348 158788 124404 285628
rect 128298 274350 128918 291922
rect 128298 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 128918 274350
rect 128298 274226 128918 274294
rect 128298 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 128918 274226
rect 128298 274102 128918 274170
rect 128298 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 128918 274102
rect 128298 273978 128918 274046
rect 128298 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 128918 273978
rect 128298 256350 128918 273922
rect 128298 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 128918 256350
rect 128298 256226 128918 256294
rect 128298 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 128918 256226
rect 128298 256102 128918 256170
rect 128298 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 128918 256102
rect 128298 255978 128918 256046
rect 128298 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 128918 255978
rect 128298 238350 128918 255922
rect 128298 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 128918 238350
rect 128298 238226 128918 238294
rect 128298 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 128918 238226
rect 128298 238102 128918 238170
rect 128298 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 128918 238102
rect 128298 237978 128918 238046
rect 128298 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 128918 237978
rect 128298 220350 128918 237922
rect 128298 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 128918 220350
rect 128298 220226 128918 220294
rect 128298 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 128918 220226
rect 128298 220102 128918 220170
rect 128298 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 128918 220102
rect 128298 219978 128918 220046
rect 128298 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 128918 219978
rect 125888 202350 126208 202384
rect 125888 202294 125958 202350
rect 126014 202294 126082 202350
rect 126138 202294 126208 202350
rect 125888 202226 126208 202294
rect 125888 202170 125958 202226
rect 126014 202170 126082 202226
rect 126138 202170 126208 202226
rect 125888 202102 126208 202170
rect 125888 202046 125958 202102
rect 126014 202046 126082 202102
rect 126138 202046 126208 202102
rect 125888 201978 126208 202046
rect 125888 201922 125958 201978
rect 126014 201922 126082 201978
rect 126138 201922 126208 201978
rect 125888 201888 126208 201922
rect 128298 202350 128918 219922
rect 132018 298350 132638 299890
rect 132018 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 132638 298350
rect 132018 298226 132638 298294
rect 132018 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 132638 298226
rect 132018 298102 132638 298170
rect 132018 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 132638 298102
rect 132018 297978 132638 298046
rect 132018 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 132638 297978
rect 132018 280350 132638 297922
rect 141248 298350 141568 298384
rect 141248 298294 141318 298350
rect 141374 298294 141442 298350
rect 141498 298294 141568 298350
rect 141248 298226 141568 298294
rect 141248 298170 141318 298226
rect 141374 298170 141442 298226
rect 141498 298170 141568 298226
rect 141248 298102 141568 298170
rect 141248 298046 141318 298102
rect 141374 298046 141442 298102
rect 141498 298046 141568 298102
rect 141248 297978 141568 298046
rect 141248 297922 141318 297978
rect 141374 297922 141442 297978
rect 141498 297922 141568 297978
rect 141248 297888 141568 297922
rect 159018 292350 159638 299890
rect 159018 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 159638 292350
rect 159018 292226 159638 292294
rect 159018 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 159638 292226
rect 159018 292102 159638 292170
rect 159018 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 159638 292102
rect 159018 291978 159638 292046
rect 159018 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 159638 291978
rect 155372 286916 155428 286926
rect 152012 286692 152068 286702
rect 149660 286580 149716 286590
rect 140252 286468 140308 286478
rect 132018 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 132638 280350
rect 132018 280226 132638 280294
rect 132018 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 132638 280226
rect 132018 280102 132638 280170
rect 132018 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 132638 280102
rect 132018 279978 132638 280046
rect 132018 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 132638 279978
rect 132018 262350 132638 279922
rect 132018 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 132638 262350
rect 132018 262226 132638 262294
rect 132018 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 132638 262226
rect 132018 262102 132638 262170
rect 132018 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 132638 262102
rect 132018 261978 132638 262046
rect 132018 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 132638 261978
rect 132018 244350 132638 261922
rect 132018 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 132638 244350
rect 132018 244226 132638 244294
rect 132018 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 132638 244226
rect 132018 244102 132638 244170
rect 132018 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 132638 244102
rect 132018 243978 132638 244046
rect 132018 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 132638 243978
rect 132018 226350 132638 243922
rect 136892 286244 136948 286254
rect 132018 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 132638 226350
rect 132018 226226 132638 226294
rect 132018 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 132638 226226
rect 132018 226102 132638 226170
rect 132018 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 132638 226102
rect 132018 225978 132638 226046
rect 132018 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 132638 225978
rect 128298 202294 128394 202350
rect 128450 202294 128518 202350
rect 128574 202294 128642 202350
rect 128698 202294 128766 202350
rect 128822 202294 128918 202350
rect 128298 202226 128918 202294
rect 128298 202170 128394 202226
rect 128450 202170 128518 202226
rect 128574 202170 128642 202226
rect 128698 202170 128766 202226
rect 128822 202170 128918 202226
rect 128298 202102 128918 202170
rect 128298 202046 128394 202102
rect 128450 202046 128518 202102
rect 128574 202046 128642 202102
rect 128698 202046 128766 202102
rect 128822 202046 128918 202102
rect 128298 201978 128918 202046
rect 128298 201922 128394 201978
rect 128450 201922 128518 201978
rect 128574 201922 128642 201978
rect 128698 201922 128766 201978
rect 128822 201922 128918 201978
rect 125888 184350 126208 184384
rect 125888 184294 125958 184350
rect 126014 184294 126082 184350
rect 126138 184294 126208 184350
rect 125888 184226 126208 184294
rect 125888 184170 125958 184226
rect 126014 184170 126082 184226
rect 126138 184170 126208 184226
rect 125888 184102 126208 184170
rect 125888 184046 125958 184102
rect 126014 184046 126082 184102
rect 126138 184046 126208 184102
rect 125888 183978 126208 184046
rect 125888 183922 125958 183978
rect 126014 183922 126082 183978
rect 126138 183922 126208 183978
rect 125888 183888 126208 183922
rect 128298 184350 128918 201922
rect 128298 184294 128394 184350
rect 128450 184294 128518 184350
rect 128574 184294 128642 184350
rect 128698 184294 128766 184350
rect 128822 184294 128918 184350
rect 128298 184226 128918 184294
rect 128298 184170 128394 184226
rect 128450 184170 128518 184226
rect 128574 184170 128642 184226
rect 128698 184170 128766 184226
rect 128822 184170 128918 184226
rect 128298 184102 128918 184170
rect 128298 184046 128394 184102
rect 128450 184046 128518 184102
rect 128574 184046 128642 184102
rect 128698 184046 128766 184102
rect 128822 184046 128918 184102
rect 128298 183978 128918 184046
rect 128298 183922 128394 183978
rect 128450 183922 128518 183978
rect 128574 183922 128642 183978
rect 128698 183922 128766 183978
rect 128822 183922 128918 183978
rect 125888 166350 126208 166384
rect 125888 166294 125958 166350
rect 126014 166294 126082 166350
rect 126138 166294 126208 166350
rect 125888 166226 126208 166294
rect 125888 166170 125958 166226
rect 126014 166170 126082 166226
rect 126138 166170 126208 166226
rect 125888 166102 126208 166170
rect 125888 166046 125958 166102
rect 126014 166046 126082 166102
rect 126138 166046 126208 166102
rect 125888 165978 126208 166046
rect 125888 165922 125958 165978
rect 126014 165922 126082 165978
rect 126138 165922 126208 165978
rect 125888 165888 126208 165922
rect 128298 166350 128918 183922
rect 128298 166294 128394 166350
rect 128450 166294 128518 166350
rect 128574 166294 128642 166350
rect 128698 166294 128766 166350
rect 128822 166294 128918 166350
rect 128298 166226 128918 166294
rect 128298 166170 128394 166226
rect 128450 166170 128518 166226
rect 128574 166170 128642 166226
rect 128698 166170 128766 166226
rect 128822 166170 128918 166226
rect 128298 166102 128918 166170
rect 128298 166046 128394 166102
rect 128450 166046 128518 166102
rect 128574 166046 128642 166102
rect 128698 166046 128766 166102
rect 128822 166046 128918 166102
rect 128298 165978 128918 166046
rect 128298 165922 128394 165978
rect 128450 165922 128518 165978
rect 128574 165922 128642 165978
rect 128698 165922 128766 165978
rect 128822 165922 128918 165978
rect 124348 158722 124404 158732
rect 121772 26002 121828 26012
rect 128298 148350 128918 165922
rect 128298 148294 128394 148350
rect 128450 148294 128518 148350
rect 128574 148294 128642 148350
rect 128698 148294 128766 148350
rect 128822 148294 128918 148350
rect 128298 148226 128918 148294
rect 128298 148170 128394 148226
rect 128450 148170 128518 148226
rect 128574 148170 128642 148226
rect 128698 148170 128766 148226
rect 128822 148170 128918 148226
rect 128298 148102 128918 148170
rect 128298 148046 128394 148102
rect 128450 148046 128518 148102
rect 128574 148046 128642 148102
rect 128698 148046 128766 148102
rect 128822 148046 128918 148102
rect 128298 147978 128918 148046
rect 128298 147922 128394 147978
rect 128450 147922 128518 147978
rect 128574 147922 128642 147978
rect 128698 147922 128766 147978
rect 128822 147922 128918 147978
rect 128298 130350 128918 147922
rect 128298 130294 128394 130350
rect 128450 130294 128518 130350
rect 128574 130294 128642 130350
rect 128698 130294 128766 130350
rect 128822 130294 128918 130350
rect 128298 130226 128918 130294
rect 128298 130170 128394 130226
rect 128450 130170 128518 130226
rect 128574 130170 128642 130226
rect 128698 130170 128766 130226
rect 128822 130170 128918 130226
rect 128298 130102 128918 130170
rect 128298 130046 128394 130102
rect 128450 130046 128518 130102
rect 128574 130046 128642 130102
rect 128698 130046 128766 130102
rect 128822 130046 128918 130102
rect 128298 129978 128918 130046
rect 128298 129922 128394 129978
rect 128450 129922 128518 129978
rect 128574 129922 128642 129978
rect 128698 129922 128766 129978
rect 128822 129922 128918 129978
rect 128298 112350 128918 129922
rect 128298 112294 128394 112350
rect 128450 112294 128518 112350
rect 128574 112294 128642 112350
rect 128698 112294 128766 112350
rect 128822 112294 128918 112350
rect 128298 112226 128918 112294
rect 128298 112170 128394 112226
rect 128450 112170 128518 112226
rect 128574 112170 128642 112226
rect 128698 112170 128766 112226
rect 128822 112170 128918 112226
rect 128298 112102 128918 112170
rect 128298 112046 128394 112102
rect 128450 112046 128518 112102
rect 128574 112046 128642 112102
rect 128698 112046 128766 112102
rect 128822 112046 128918 112102
rect 128298 111978 128918 112046
rect 128298 111922 128394 111978
rect 128450 111922 128518 111978
rect 128574 111922 128642 111978
rect 128698 111922 128766 111978
rect 128822 111922 128918 111978
rect 128298 94350 128918 111922
rect 128298 94294 128394 94350
rect 128450 94294 128518 94350
rect 128574 94294 128642 94350
rect 128698 94294 128766 94350
rect 128822 94294 128918 94350
rect 128298 94226 128918 94294
rect 128298 94170 128394 94226
rect 128450 94170 128518 94226
rect 128574 94170 128642 94226
rect 128698 94170 128766 94226
rect 128822 94170 128918 94226
rect 128298 94102 128918 94170
rect 128298 94046 128394 94102
rect 128450 94046 128518 94102
rect 128574 94046 128642 94102
rect 128698 94046 128766 94102
rect 128822 94046 128918 94102
rect 128298 93978 128918 94046
rect 128298 93922 128394 93978
rect 128450 93922 128518 93978
rect 128574 93922 128642 93978
rect 128698 93922 128766 93978
rect 128822 93922 128918 93978
rect 128298 76350 128918 93922
rect 128298 76294 128394 76350
rect 128450 76294 128518 76350
rect 128574 76294 128642 76350
rect 128698 76294 128766 76350
rect 128822 76294 128918 76350
rect 128298 76226 128918 76294
rect 128298 76170 128394 76226
rect 128450 76170 128518 76226
rect 128574 76170 128642 76226
rect 128698 76170 128766 76226
rect 128822 76170 128918 76226
rect 128298 76102 128918 76170
rect 128298 76046 128394 76102
rect 128450 76046 128518 76102
rect 128574 76046 128642 76102
rect 128698 76046 128766 76102
rect 128822 76046 128918 76102
rect 128298 75978 128918 76046
rect 128298 75922 128394 75978
rect 128450 75922 128518 75978
rect 128574 75922 128642 75978
rect 128698 75922 128766 75978
rect 128822 75922 128918 75978
rect 128298 58350 128918 75922
rect 128298 58294 128394 58350
rect 128450 58294 128518 58350
rect 128574 58294 128642 58350
rect 128698 58294 128766 58350
rect 128822 58294 128918 58350
rect 128298 58226 128918 58294
rect 128298 58170 128394 58226
rect 128450 58170 128518 58226
rect 128574 58170 128642 58226
rect 128698 58170 128766 58226
rect 128822 58170 128918 58226
rect 128298 58102 128918 58170
rect 128298 58046 128394 58102
rect 128450 58046 128518 58102
rect 128574 58046 128642 58102
rect 128698 58046 128766 58102
rect 128822 58046 128918 58102
rect 128298 57978 128918 58046
rect 128298 57922 128394 57978
rect 128450 57922 128518 57978
rect 128574 57922 128642 57978
rect 128698 57922 128766 57978
rect 128822 57922 128918 57978
rect 128298 40350 128918 57922
rect 128298 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 128918 40350
rect 128298 40226 128918 40294
rect 128298 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 128918 40226
rect 128298 40102 128918 40170
rect 128298 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 128918 40102
rect 128298 39978 128918 40046
rect 128298 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 128918 39978
rect 119196 4162 119252 4172
rect 128298 22350 128918 39922
rect 128298 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 128918 22350
rect 128298 22226 128918 22294
rect 128298 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 128918 22226
rect 128298 22102 128918 22170
rect 128298 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 128918 22102
rect 128298 21978 128918 22046
rect 128298 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 128918 21978
rect 128298 4350 128918 21922
rect 130172 212772 130228 212782
rect 130172 4676 130228 212716
rect 132018 208350 132638 225922
rect 132018 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 132638 208350
rect 132018 208226 132638 208294
rect 132018 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 132638 208226
rect 132018 208102 132638 208170
rect 132018 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 132638 208102
rect 132018 207978 132638 208046
rect 132018 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 132638 207978
rect 132018 190350 132638 207922
rect 132018 190294 132114 190350
rect 132170 190294 132238 190350
rect 132294 190294 132362 190350
rect 132418 190294 132486 190350
rect 132542 190294 132638 190350
rect 132018 190226 132638 190294
rect 132018 190170 132114 190226
rect 132170 190170 132238 190226
rect 132294 190170 132362 190226
rect 132418 190170 132486 190226
rect 132542 190170 132638 190226
rect 132018 190102 132638 190170
rect 132018 190046 132114 190102
rect 132170 190046 132238 190102
rect 132294 190046 132362 190102
rect 132418 190046 132486 190102
rect 132542 190046 132638 190102
rect 132018 189978 132638 190046
rect 132018 189922 132114 189978
rect 132170 189922 132238 189978
rect 132294 189922 132362 189978
rect 132418 189922 132486 189978
rect 132542 189922 132638 189978
rect 132018 172350 132638 189922
rect 132018 172294 132114 172350
rect 132170 172294 132238 172350
rect 132294 172294 132362 172350
rect 132418 172294 132486 172350
rect 132542 172294 132638 172350
rect 132018 172226 132638 172294
rect 132018 172170 132114 172226
rect 132170 172170 132238 172226
rect 132294 172170 132362 172226
rect 132418 172170 132486 172226
rect 132542 172170 132638 172226
rect 132018 172102 132638 172170
rect 132018 172046 132114 172102
rect 132170 172046 132238 172102
rect 132294 172046 132362 172102
rect 132418 172046 132486 172102
rect 132542 172046 132638 172102
rect 132018 171978 132638 172046
rect 132018 171922 132114 171978
rect 132170 171922 132238 171978
rect 132294 171922 132362 171978
rect 132418 171922 132486 171978
rect 132542 171922 132638 171978
rect 132018 154350 132638 171922
rect 132018 154294 132114 154350
rect 132170 154294 132238 154350
rect 132294 154294 132362 154350
rect 132418 154294 132486 154350
rect 132542 154294 132638 154350
rect 132018 154226 132638 154294
rect 132018 154170 132114 154226
rect 132170 154170 132238 154226
rect 132294 154170 132362 154226
rect 132418 154170 132486 154226
rect 132542 154170 132638 154226
rect 132018 154102 132638 154170
rect 132018 154046 132114 154102
rect 132170 154046 132238 154102
rect 132294 154046 132362 154102
rect 132418 154046 132486 154102
rect 132542 154046 132638 154102
rect 132018 153978 132638 154046
rect 132018 153922 132114 153978
rect 132170 153922 132238 153978
rect 132294 153922 132362 153978
rect 132418 153922 132486 153978
rect 132542 153922 132638 153978
rect 130956 142324 131012 142356
rect 130956 142252 131012 142262
rect 130172 4610 130228 4620
rect 132018 136350 132638 153922
rect 132018 136294 132114 136350
rect 132170 136294 132238 136350
rect 132294 136294 132362 136350
rect 132418 136294 132486 136350
rect 132542 136294 132638 136350
rect 132018 136226 132638 136294
rect 132018 136170 132114 136226
rect 132170 136170 132238 136226
rect 132294 136170 132362 136226
rect 132418 136170 132486 136226
rect 132542 136170 132638 136226
rect 132018 136102 132638 136170
rect 132018 136046 132114 136102
rect 132170 136046 132238 136102
rect 132294 136046 132362 136102
rect 132418 136046 132486 136102
rect 132542 136046 132638 136102
rect 132018 135978 132638 136046
rect 132018 135922 132114 135978
rect 132170 135922 132238 135978
rect 132294 135922 132362 135978
rect 132418 135922 132486 135978
rect 132542 135922 132638 135978
rect 132018 118350 132638 135922
rect 132018 118294 132114 118350
rect 132170 118294 132238 118350
rect 132294 118294 132362 118350
rect 132418 118294 132486 118350
rect 132542 118294 132638 118350
rect 132018 118226 132638 118294
rect 132018 118170 132114 118226
rect 132170 118170 132238 118226
rect 132294 118170 132362 118226
rect 132418 118170 132486 118226
rect 132542 118170 132638 118226
rect 132018 118102 132638 118170
rect 132018 118046 132114 118102
rect 132170 118046 132238 118102
rect 132294 118046 132362 118102
rect 132418 118046 132486 118102
rect 132542 118046 132638 118102
rect 132018 117978 132638 118046
rect 132018 117922 132114 117978
rect 132170 117922 132238 117978
rect 132294 117922 132362 117978
rect 132418 117922 132486 117978
rect 132542 117922 132638 117978
rect 132018 100350 132638 117922
rect 132018 100294 132114 100350
rect 132170 100294 132238 100350
rect 132294 100294 132362 100350
rect 132418 100294 132486 100350
rect 132542 100294 132638 100350
rect 132018 100226 132638 100294
rect 132018 100170 132114 100226
rect 132170 100170 132238 100226
rect 132294 100170 132362 100226
rect 132418 100170 132486 100226
rect 132542 100170 132638 100226
rect 132018 100102 132638 100170
rect 132018 100046 132114 100102
rect 132170 100046 132238 100102
rect 132294 100046 132362 100102
rect 132418 100046 132486 100102
rect 132542 100046 132638 100102
rect 132018 99978 132638 100046
rect 132018 99922 132114 99978
rect 132170 99922 132238 99978
rect 132294 99922 132362 99978
rect 132418 99922 132486 99978
rect 132542 99922 132638 99978
rect 132018 82350 132638 99922
rect 132018 82294 132114 82350
rect 132170 82294 132238 82350
rect 132294 82294 132362 82350
rect 132418 82294 132486 82350
rect 132542 82294 132638 82350
rect 132018 82226 132638 82294
rect 132018 82170 132114 82226
rect 132170 82170 132238 82226
rect 132294 82170 132362 82226
rect 132418 82170 132486 82226
rect 132542 82170 132638 82226
rect 132018 82102 132638 82170
rect 132018 82046 132114 82102
rect 132170 82046 132238 82102
rect 132294 82046 132362 82102
rect 132418 82046 132486 82102
rect 132542 82046 132638 82102
rect 132018 81978 132638 82046
rect 132018 81922 132114 81978
rect 132170 81922 132238 81978
rect 132294 81922 132362 81978
rect 132418 81922 132486 81978
rect 132542 81922 132638 81978
rect 132018 64350 132638 81922
rect 132018 64294 132114 64350
rect 132170 64294 132238 64350
rect 132294 64294 132362 64350
rect 132418 64294 132486 64350
rect 132542 64294 132638 64350
rect 132018 64226 132638 64294
rect 132018 64170 132114 64226
rect 132170 64170 132238 64226
rect 132294 64170 132362 64226
rect 132418 64170 132486 64226
rect 132542 64170 132638 64226
rect 132018 64102 132638 64170
rect 132018 64046 132114 64102
rect 132170 64046 132238 64102
rect 132294 64046 132362 64102
rect 132418 64046 132486 64102
rect 132542 64046 132638 64102
rect 132018 63978 132638 64046
rect 132018 63922 132114 63978
rect 132170 63922 132238 63978
rect 132294 63922 132362 63978
rect 132418 63922 132486 63978
rect 132542 63922 132638 63978
rect 132018 46350 132638 63922
rect 132018 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 132638 46350
rect 132018 46226 132638 46294
rect 132018 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 132638 46226
rect 132018 46102 132638 46170
rect 132018 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 132638 46102
rect 132018 45978 132638 46046
rect 132018 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 132638 45978
rect 132018 28350 132638 45922
rect 132018 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 132638 28350
rect 132018 28226 132638 28294
rect 132018 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 132638 28226
rect 132018 28102 132638 28170
rect 132018 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 132638 28102
rect 132018 27978 132638 28046
rect 132018 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 132638 27978
rect 132018 10350 132638 27922
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 -1120 132638 9922
rect 133532 231028 133588 231038
rect 133532 4004 133588 230972
rect 135212 210980 135268 210990
rect 135212 4116 135268 210924
rect 136892 6020 136948 286188
rect 138572 285684 138628 285694
rect 138572 15988 138628 285628
rect 138572 15922 138628 15932
rect 136892 5954 136948 5964
rect 140252 5124 140308 286412
rect 147980 286356 148036 286366
rect 147868 285684 147924 285694
rect 141248 190350 141568 190384
rect 141248 190294 141318 190350
rect 141374 190294 141442 190350
rect 141498 190294 141568 190350
rect 141248 190226 141568 190294
rect 141248 190170 141318 190226
rect 141374 190170 141442 190226
rect 141498 190170 141568 190226
rect 141248 190102 141568 190170
rect 141248 190046 141318 190102
rect 141374 190046 141442 190102
rect 141498 190046 141568 190102
rect 141248 189978 141568 190046
rect 141248 189922 141318 189978
rect 141374 189922 141442 189978
rect 141498 189922 141568 189978
rect 141248 189888 141568 189922
rect 141248 172350 141568 172384
rect 141248 172294 141318 172350
rect 141374 172294 141442 172350
rect 141498 172294 141568 172350
rect 141248 172226 141568 172294
rect 141248 172170 141318 172226
rect 141374 172170 141442 172226
rect 141498 172170 141568 172226
rect 141248 172102 141568 172170
rect 141248 172046 141318 172102
rect 141374 172046 141442 172102
rect 141498 172046 141568 172102
rect 141248 171978 141568 172046
rect 141248 171922 141318 171978
rect 141374 171922 141442 171978
rect 141498 171922 141568 171978
rect 141248 171888 141568 171922
rect 144508 155540 144564 155550
rect 144508 142436 144564 155484
rect 144732 152180 144788 152190
rect 144732 142772 144788 152124
rect 144732 142678 144788 142716
rect 144732 142612 144788 142622
rect 144508 142370 144564 142380
rect 145404 141204 145460 141214
rect 145404 140878 145460 141148
rect 145404 140812 145460 140822
rect 145788 130350 146264 130384
rect 145788 130294 145812 130350
rect 145868 130294 145936 130350
rect 145992 130294 146060 130350
rect 146116 130294 146184 130350
rect 146240 130294 146264 130350
rect 145788 130226 146264 130294
rect 145788 130170 145812 130226
rect 145868 130170 145936 130226
rect 145992 130170 146060 130226
rect 146116 130170 146184 130226
rect 146240 130170 146264 130226
rect 145788 130102 146264 130170
rect 145788 130046 145812 130102
rect 145868 130046 145936 130102
rect 145992 130046 146060 130102
rect 146116 130046 146184 130102
rect 146240 130046 146264 130102
rect 145788 129978 146264 130046
rect 145788 129922 145812 129978
rect 145868 129922 145936 129978
rect 145992 129922 146060 129978
rect 146116 129922 146184 129978
rect 146240 129922 146264 129978
rect 145788 129888 146264 129922
rect 146588 118350 147064 118384
rect 146588 118294 146612 118350
rect 146668 118294 146736 118350
rect 146792 118294 146860 118350
rect 146916 118294 146984 118350
rect 147040 118294 147064 118350
rect 146588 118226 147064 118294
rect 146588 118170 146612 118226
rect 146668 118170 146736 118226
rect 146792 118170 146860 118226
rect 146916 118170 146984 118226
rect 147040 118170 147064 118226
rect 146588 118102 147064 118170
rect 146588 118046 146612 118102
rect 146668 118046 146736 118102
rect 146792 118046 146860 118102
rect 146916 118046 146984 118102
rect 147040 118046 147064 118102
rect 146588 117978 147064 118046
rect 146588 117922 146612 117978
rect 146668 117922 146736 117978
rect 146792 117922 146860 117978
rect 146916 117922 146984 117978
rect 147040 117922 147064 117978
rect 146588 117888 147064 117922
rect 145788 112350 146264 112384
rect 145788 112294 145812 112350
rect 145868 112294 145936 112350
rect 145992 112294 146060 112350
rect 146116 112294 146184 112350
rect 146240 112294 146264 112350
rect 145788 112226 146264 112294
rect 145788 112170 145812 112226
rect 145868 112170 145936 112226
rect 145992 112170 146060 112226
rect 146116 112170 146184 112226
rect 146240 112170 146264 112226
rect 145788 112102 146264 112170
rect 145788 112046 145812 112102
rect 145868 112046 145936 112102
rect 145992 112046 146060 112102
rect 146116 112046 146184 112102
rect 146240 112046 146264 112102
rect 145788 111978 146264 112046
rect 145788 111922 145812 111978
rect 145868 111922 145936 111978
rect 145992 111922 146060 111978
rect 146116 111922 146184 111978
rect 146240 111922 146264 111978
rect 145788 111888 146264 111922
rect 146588 100350 147064 100384
rect 146588 100294 146612 100350
rect 146668 100294 146736 100350
rect 146792 100294 146860 100350
rect 146916 100294 146984 100350
rect 147040 100294 147064 100350
rect 146588 100226 147064 100294
rect 146588 100170 146612 100226
rect 146668 100170 146736 100226
rect 146792 100170 146860 100226
rect 146916 100170 146984 100226
rect 147040 100170 147064 100226
rect 146588 100102 147064 100170
rect 146588 100046 146612 100102
rect 146668 100046 146736 100102
rect 146792 100046 146860 100102
rect 146916 100046 146984 100102
rect 147040 100046 147064 100102
rect 146588 99978 147064 100046
rect 146588 99922 146612 99978
rect 146668 99922 146736 99978
rect 146792 99922 146860 99978
rect 146916 99922 146984 99978
rect 147040 99922 147064 99978
rect 146588 99888 147064 99922
rect 145788 94350 146264 94384
rect 145788 94294 145812 94350
rect 145868 94294 145936 94350
rect 145992 94294 146060 94350
rect 146116 94294 146184 94350
rect 146240 94294 146264 94350
rect 145788 94226 146264 94294
rect 145788 94170 145812 94226
rect 145868 94170 145936 94226
rect 145992 94170 146060 94226
rect 146116 94170 146184 94226
rect 146240 94170 146264 94226
rect 145788 94102 146264 94170
rect 145788 94046 145812 94102
rect 145868 94046 145936 94102
rect 145992 94046 146060 94102
rect 146116 94046 146184 94102
rect 146240 94046 146264 94102
rect 145788 93978 146264 94046
rect 145788 93922 145812 93978
rect 145868 93922 145936 93978
rect 145992 93922 146060 93978
rect 146116 93922 146184 93978
rect 146240 93922 146264 93978
rect 145788 93888 146264 93922
rect 146588 82350 147064 82384
rect 146588 82294 146612 82350
rect 146668 82294 146736 82350
rect 146792 82294 146860 82350
rect 146916 82294 146984 82350
rect 147040 82294 147064 82350
rect 146588 82226 147064 82294
rect 146588 82170 146612 82226
rect 146668 82170 146736 82226
rect 146792 82170 146860 82226
rect 146916 82170 146984 82226
rect 147040 82170 147064 82226
rect 146588 82102 147064 82170
rect 146588 82046 146612 82102
rect 146668 82046 146736 82102
rect 146792 82046 146860 82102
rect 146916 82046 146984 82102
rect 147040 82046 147064 82102
rect 146588 81978 147064 82046
rect 146588 81922 146612 81978
rect 146668 81922 146736 81978
rect 146792 81922 146860 81978
rect 146916 81922 146984 81978
rect 147040 81922 147064 81978
rect 146588 81888 147064 81922
rect 145788 76350 146264 76384
rect 145788 76294 145812 76350
rect 145868 76294 145936 76350
rect 145992 76294 146060 76350
rect 146116 76294 146184 76350
rect 146240 76294 146264 76350
rect 145788 76226 146264 76294
rect 145788 76170 145812 76226
rect 145868 76170 145936 76226
rect 145992 76170 146060 76226
rect 146116 76170 146184 76226
rect 146240 76170 146264 76226
rect 145788 76102 146264 76170
rect 145788 76046 145812 76102
rect 145868 76046 145936 76102
rect 145992 76046 146060 76102
rect 146116 76046 146184 76102
rect 146240 76046 146264 76102
rect 145788 75978 146264 76046
rect 145788 75922 145812 75978
rect 145868 75922 145936 75978
rect 145992 75922 146060 75978
rect 146116 75922 146184 75978
rect 146240 75922 146264 75978
rect 145788 75888 146264 75922
rect 146588 64350 147064 64384
rect 146588 64294 146612 64350
rect 146668 64294 146736 64350
rect 146792 64294 146860 64350
rect 146916 64294 146984 64350
rect 147040 64294 147064 64350
rect 146588 64226 147064 64294
rect 146588 64170 146612 64226
rect 146668 64170 146736 64226
rect 146792 64170 146860 64226
rect 146916 64170 146984 64226
rect 147040 64170 147064 64226
rect 146588 64102 147064 64170
rect 146588 64046 146612 64102
rect 146668 64046 146736 64102
rect 146792 64046 146860 64102
rect 146916 64046 146984 64102
rect 147040 64046 147064 64102
rect 146588 63978 147064 64046
rect 146588 63922 146612 63978
rect 146668 63922 146736 63978
rect 146792 63922 146860 63978
rect 146916 63922 146984 63978
rect 147040 63922 147064 63978
rect 146588 63888 147064 63922
rect 145788 58350 146264 58384
rect 145788 58294 145812 58350
rect 145868 58294 145936 58350
rect 145992 58294 146060 58350
rect 146116 58294 146184 58350
rect 146240 58294 146264 58350
rect 145788 58226 146264 58294
rect 145788 58170 145812 58226
rect 145868 58170 145936 58226
rect 145992 58170 146060 58226
rect 146116 58170 146184 58226
rect 146240 58170 146264 58226
rect 145788 58102 146264 58170
rect 145788 58046 145812 58102
rect 145868 58046 145936 58102
rect 145992 58046 146060 58102
rect 146116 58046 146184 58102
rect 146240 58046 146264 58102
rect 145788 57978 146264 58046
rect 145788 57922 145812 57978
rect 145868 57922 145936 57978
rect 145992 57922 146060 57978
rect 146116 57922 146184 57978
rect 146240 57922 146264 57978
rect 145788 57888 146264 57922
rect 146588 46350 147064 46384
rect 146588 46294 146612 46350
rect 146668 46294 146736 46350
rect 146792 46294 146860 46350
rect 146916 46294 146984 46350
rect 147040 46294 147064 46350
rect 146588 46226 147064 46294
rect 146588 46170 146612 46226
rect 146668 46170 146736 46226
rect 146792 46170 146860 46226
rect 146916 46170 146984 46226
rect 147040 46170 147064 46226
rect 146588 46102 147064 46170
rect 146588 46046 146612 46102
rect 146668 46046 146736 46102
rect 146792 46046 146860 46102
rect 146916 46046 146984 46102
rect 147040 46046 147064 46102
rect 146588 45978 147064 46046
rect 146588 45922 146612 45978
rect 146668 45922 146736 45978
rect 146792 45922 146860 45978
rect 146916 45922 146984 45978
rect 147040 45922 147064 45978
rect 146588 45888 147064 45922
rect 147868 7588 147924 285628
rect 147980 24388 148036 286300
rect 147980 24322 148036 24332
rect 149548 286244 149604 286254
rect 149548 7700 149604 286188
rect 149660 36148 149716 286524
rect 149772 286020 149828 286030
rect 149772 39508 149828 285964
rect 152012 40292 152068 286636
rect 152908 285796 152964 285806
rect 152012 40226 152068 40236
rect 152124 167338 152180 167348
rect 149772 39442 149828 39452
rect 149660 36082 149716 36092
rect 149548 7634 149604 7644
rect 147868 7522 147924 7532
rect 140252 5058 140308 5068
rect 152124 5012 152180 167282
rect 152908 5908 152964 285740
rect 153020 285684 153076 285694
rect 153020 12628 153076 285628
rect 154588 285684 154644 285694
rect 154588 37940 154644 285628
rect 154588 37874 154644 37884
rect 155372 36260 155428 286860
rect 159018 274350 159638 291922
rect 162738 298350 163358 299890
rect 162738 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 163358 298350
rect 162738 298226 163358 298294
rect 162738 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 163358 298226
rect 162738 298102 163358 298170
rect 162738 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 163358 298102
rect 162738 297978 163358 298046
rect 162738 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 163358 297978
rect 159018 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 159638 274350
rect 159018 274226 159638 274294
rect 159018 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 159638 274226
rect 159018 274102 159638 274170
rect 159018 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 159638 274102
rect 159018 273978 159638 274046
rect 159018 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 159638 273978
rect 159018 256350 159638 273922
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 156608 202350 156928 202384
rect 156608 202294 156678 202350
rect 156734 202294 156802 202350
rect 156858 202294 156928 202350
rect 156608 202226 156928 202294
rect 156608 202170 156678 202226
rect 156734 202170 156802 202226
rect 156858 202170 156928 202226
rect 156608 202102 156928 202170
rect 156608 202046 156678 202102
rect 156734 202046 156802 202102
rect 156858 202046 156928 202102
rect 156608 201978 156928 202046
rect 156608 201922 156678 201978
rect 156734 201922 156802 201978
rect 156858 201922 156928 201978
rect 156608 201888 156928 201922
rect 159018 202350 159638 219922
rect 159018 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 159638 202350
rect 159018 202226 159638 202294
rect 159018 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 159638 202226
rect 159018 202102 159638 202170
rect 159018 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 159638 202102
rect 159018 201978 159638 202046
rect 159018 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 159638 201978
rect 156608 184350 156928 184384
rect 156608 184294 156678 184350
rect 156734 184294 156802 184350
rect 156858 184294 156928 184350
rect 156608 184226 156928 184294
rect 156608 184170 156678 184226
rect 156734 184170 156802 184226
rect 156858 184170 156928 184226
rect 156608 184102 156928 184170
rect 156608 184046 156678 184102
rect 156734 184046 156802 184102
rect 156858 184046 156928 184102
rect 156608 183978 156928 184046
rect 156608 183922 156678 183978
rect 156734 183922 156802 183978
rect 156858 183922 156928 183978
rect 156608 183888 156928 183922
rect 159018 184350 159638 201922
rect 159018 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 159638 184350
rect 159018 184226 159638 184294
rect 159018 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 159638 184226
rect 159018 184102 159638 184170
rect 159018 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 159638 184102
rect 159018 183978 159638 184046
rect 159018 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 159638 183978
rect 157052 168778 157108 168788
rect 156608 166350 156928 166384
rect 156608 166294 156678 166350
rect 156734 166294 156802 166350
rect 156858 166294 156928 166350
rect 156608 166226 156928 166294
rect 156608 166170 156678 166226
rect 156734 166170 156802 166226
rect 156858 166170 156928 166226
rect 156608 166102 156928 166170
rect 156608 166046 156678 166102
rect 156734 166046 156802 166102
rect 156858 166046 156928 166102
rect 156608 165978 156928 166046
rect 156608 165922 156678 165978
rect 156734 165922 156802 165978
rect 156858 165922 156928 165978
rect 156608 165888 156928 165922
rect 155372 36194 155428 36204
rect 155484 150612 155540 150622
rect 153020 12562 153076 12572
rect 152908 5842 152964 5852
rect 135212 4050 135268 4060
rect 137228 4978 137284 4988
rect 152124 4946 152180 4956
rect 155484 4978 155540 150556
rect 133532 3938 133588 3948
rect 137228 3444 137284 4922
rect 155484 4912 155540 4922
rect 143612 4788 143668 4798
rect 143612 4116 143668 4732
rect 157052 4228 157108 168722
rect 157052 4162 157108 4172
rect 159018 166350 159638 183922
rect 159018 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 159638 166350
rect 159018 166226 159638 166294
rect 159018 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 159638 166226
rect 159018 166102 159638 166170
rect 159018 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 159638 166102
rect 159018 165978 159638 166046
rect 159018 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 159638 165978
rect 159018 148350 159638 165922
rect 159018 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 159638 148350
rect 159018 148226 159638 148294
rect 159018 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 159638 148226
rect 159018 148102 159638 148170
rect 159018 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 159638 148102
rect 159018 147978 159638 148046
rect 159018 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 159638 147978
rect 159018 130350 159638 147922
rect 159018 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 159638 130350
rect 159018 130226 159638 130294
rect 159018 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 159638 130226
rect 159018 130102 159638 130170
rect 159018 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 159638 130102
rect 159018 129978 159638 130046
rect 159018 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 159638 129978
rect 159018 112350 159638 129922
rect 159018 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 159638 112350
rect 159018 112226 159638 112294
rect 159018 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 159638 112226
rect 159018 112102 159638 112170
rect 159018 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 159638 112102
rect 159018 111978 159638 112046
rect 159018 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 159638 111978
rect 159018 94350 159638 111922
rect 159018 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 159638 94350
rect 159018 94226 159638 94294
rect 159018 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 159638 94226
rect 159018 94102 159638 94170
rect 159018 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 159638 94102
rect 159018 93978 159638 94046
rect 159018 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 159638 93978
rect 159018 76350 159638 93922
rect 159018 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 159638 76350
rect 159018 76226 159638 76294
rect 159018 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 159638 76226
rect 159018 76102 159638 76170
rect 159018 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 159638 76102
rect 159018 75978 159638 76046
rect 159018 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 159638 75978
rect 159018 58350 159638 75922
rect 159018 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 159638 58350
rect 159018 58226 159638 58294
rect 159018 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 159638 58226
rect 159018 58102 159638 58170
rect 159018 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 159638 58102
rect 159018 57978 159638 58046
rect 159018 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 159638 57978
rect 159018 40350 159638 57922
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 159018 22350 159638 39922
rect 159740 285684 159796 285694
rect 159740 37828 159796 285628
rect 162738 280350 163358 297922
rect 171968 298350 172288 298384
rect 171968 298294 172038 298350
rect 172094 298294 172162 298350
rect 172218 298294 172288 298350
rect 171968 298226 172288 298294
rect 171968 298170 172038 298226
rect 172094 298170 172162 298226
rect 172218 298170 172288 298226
rect 171968 298102 172288 298170
rect 171968 298046 172038 298102
rect 172094 298046 172162 298102
rect 172218 298046 172288 298102
rect 171968 297978 172288 298046
rect 171968 297922 172038 297978
rect 172094 297922 172162 297978
rect 172218 297922 172288 297978
rect 171968 297888 172288 297922
rect 189738 292350 190358 299890
rect 189738 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 190358 292350
rect 189738 292226 190358 292294
rect 189738 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 190358 292226
rect 189738 292102 190358 292170
rect 189738 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 190358 292102
rect 189738 291978 190358 292046
rect 189738 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 190358 291978
rect 180572 287028 180628 287038
rect 177212 286916 177268 286926
rect 167132 286804 167188 286814
rect 162738 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 163358 280350
rect 162738 280226 163358 280294
rect 162738 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 163358 280226
rect 162738 280102 163358 280170
rect 162738 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 163358 280102
rect 162738 279978 163358 280046
rect 162738 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 163358 279978
rect 162738 262350 163358 279922
rect 162738 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 163358 262350
rect 162738 262226 163358 262294
rect 162738 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 163358 262226
rect 162738 262102 163358 262170
rect 162738 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 163358 262102
rect 162738 261978 163358 262046
rect 162738 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 163358 261978
rect 162738 244350 163358 261922
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162738 226350 163358 243922
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 162738 208350 163358 225922
rect 162738 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 163358 208350
rect 162738 208226 163358 208294
rect 162738 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 163358 208226
rect 162738 208102 163358 208170
rect 162738 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 163358 208102
rect 162738 207978 163358 208046
rect 162738 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 163358 207978
rect 162738 190350 163358 207922
rect 162738 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 163358 190350
rect 162738 190226 163358 190294
rect 162738 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 163358 190226
rect 162738 190102 163358 190170
rect 162738 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 163358 190102
rect 162738 189978 163358 190046
rect 162738 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 163358 189978
rect 159740 37762 159796 37772
rect 160412 173818 160468 173828
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 159018 4350 159638 21922
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 160412 4340 160468 173762
rect 162738 172350 163358 189922
rect 162738 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 163358 172350
rect 162738 172226 163358 172294
rect 162738 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 163358 172226
rect 162738 172102 163358 172170
rect 162738 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 163358 172102
rect 162738 171978 163358 172046
rect 162738 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 163358 171978
rect 162738 154350 163358 171922
rect 162738 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 163358 154350
rect 162738 154226 163358 154294
rect 162738 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 163358 154226
rect 162738 154102 163358 154170
rect 162738 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 163358 154102
rect 162738 153978 163358 154046
rect 162738 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 163358 153978
rect 162738 136350 163358 153922
rect 164668 285684 164724 285694
rect 164668 147140 164724 285628
rect 164668 147074 164724 147084
rect 167132 144228 167188 286748
rect 168812 286580 168868 286590
rect 167132 144162 167188 144172
rect 167916 170578 167972 170588
rect 164444 142138 164500 142148
rect 164444 141316 164500 142082
rect 164444 141250 164500 141260
rect 162738 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 163358 136350
rect 162738 136226 163358 136294
rect 162738 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 163358 136226
rect 162738 136102 163358 136170
rect 162738 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 163358 136102
rect 162738 135978 163358 136046
rect 162738 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 163358 135978
rect 161106 130350 161582 130384
rect 161106 130294 161130 130350
rect 161186 130294 161254 130350
rect 161310 130294 161378 130350
rect 161434 130294 161502 130350
rect 161558 130294 161582 130350
rect 161106 130226 161582 130294
rect 161106 130170 161130 130226
rect 161186 130170 161254 130226
rect 161310 130170 161378 130226
rect 161434 130170 161502 130226
rect 161558 130170 161582 130226
rect 161106 130102 161582 130170
rect 161106 130046 161130 130102
rect 161186 130046 161254 130102
rect 161310 130046 161378 130102
rect 161434 130046 161502 130102
rect 161558 130046 161582 130102
rect 161106 129978 161582 130046
rect 161106 129922 161130 129978
rect 161186 129922 161254 129978
rect 161310 129922 161378 129978
rect 161434 129922 161502 129978
rect 161558 129922 161582 129978
rect 161106 129888 161582 129922
rect 161906 118350 162382 118384
rect 161906 118294 161930 118350
rect 161986 118294 162054 118350
rect 162110 118294 162178 118350
rect 162234 118294 162302 118350
rect 162358 118294 162382 118350
rect 161906 118226 162382 118294
rect 161906 118170 161930 118226
rect 161986 118170 162054 118226
rect 162110 118170 162178 118226
rect 162234 118170 162302 118226
rect 162358 118170 162382 118226
rect 161906 118102 162382 118170
rect 161906 118046 161930 118102
rect 161986 118046 162054 118102
rect 162110 118046 162178 118102
rect 162234 118046 162302 118102
rect 162358 118046 162382 118102
rect 161906 117978 162382 118046
rect 161906 117922 161930 117978
rect 161986 117922 162054 117978
rect 162110 117922 162178 117978
rect 162234 117922 162302 117978
rect 162358 117922 162382 117978
rect 161906 117888 162382 117922
rect 162738 118350 163358 135922
rect 162738 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 163358 118350
rect 162738 118226 163358 118294
rect 162738 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 163358 118226
rect 162738 118102 163358 118170
rect 162738 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 163358 118102
rect 162738 117978 163358 118046
rect 162738 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 163358 117978
rect 161106 112350 161582 112384
rect 161106 112294 161130 112350
rect 161186 112294 161254 112350
rect 161310 112294 161378 112350
rect 161434 112294 161502 112350
rect 161558 112294 161582 112350
rect 161106 112226 161582 112294
rect 161106 112170 161130 112226
rect 161186 112170 161254 112226
rect 161310 112170 161378 112226
rect 161434 112170 161502 112226
rect 161558 112170 161582 112226
rect 161106 112102 161582 112170
rect 161106 112046 161130 112102
rect 161186 112046 161254 112102
rect 161310 112046 161378 112102
rect 161434 112046 161502 112102
rect 161558 112046 161582 112102
rect 161106 111978 161582 112046
rect 161106 111922 161130 111978
rect 161186 111922 161254 111978
rect 161310 111922 161378 111978
rect 161434 111922 161502 111978
rect 161558 111922 161582 111978
rect 161106 111888 161582 111922
rect 161906 100350 162382 100384
rect 161906 100294 161930 100350
rect 161986 100294 162054 100350
rect 162110 100294 162178 100350
rect 162234 100294 162302 100350
rect 162358 100294 162382 100350
rect 161906 100226 162382 100294
rect 161906 100170 161930 100226
rect 161986 100170 162054 100226
rect 162110 100170 162178 100226
rect 162234 100170 162302 100226
rect 162358 100170 162382 100226
rect 161906 100102 162382 100170
rect 161906 100046 161930 100102
rect 161986 100046 162054 100102
rect 162110 100046 162178 100102
rect 162234 100046 162302 100102
rect 162358 100046 162382 100102
rect 161906 99978 162382 100046
rect 161906 99922 161930 99978
rect 161986 99922 162054 99978
rect 162110 99922 162178 99978
rect 162234 99922 162302 99978
rect 162358 99922 162382 99978
rect 161906 99888 162382 99922
rect 162738 100350 163358 117922
rect 162738 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 163358 100350
rect 162738 100226 163358 100294
rect 162738 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 163358 100226
rect 162738 100102 163358 100170
rect 162738 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 163358 100102
rect 162738 99978 163358 100046
rect 162738 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 163358 99978
rect 161106 94350 161582 94384
rect 161106 94294 161130 94350
rect 161186 94294 161254 94350
rect 161310 94294 161378 94350
rect 161434 94294 161502 94350
rect 161558 94294 161582 94350
rect 161106 94226 161582 94294
rect 161106 94170 161130 94226
rect 161186 94170 161254 94226
rect 161310 94170 161378 94226
rect 161434 94170 161502 94226
rect 161558 94170 161582 94226
rect 161106 94102 161582 94170
rect 161106 94046 161130 94102
rect 161186 94046 161254 94102
rect 161310 94046 161378 94102
rect 161434 94046 161502 94102
rect 161558 94046 161582 94102
rect 161106 93978 161582 94046
rect 161106 93922 161130 93978
rect 161186 93922 161254 93978
rect 161310 93922 161378 93978
rect 161434 93922 161502 93978
rect 161558 93922 161582 93978
rect 161106 93888 161582 93922
rect 161906 82350 162382 82384
rect 161906 82294 161930 82350
rect 161986 82294 162054 82350
rect 162110 82294 162178 82350
rect 162234 82294 162302 82350
rect 162358 82294 162382 82350
rect 161906 82226 162382 82294
rect 161906 82170 161930 82226
rect 161986 82170 162054 82226
rect 162110 82170 162178 82226
rect 162234 82170 162302 82226
rect 162358 82170 162382 82226
rect 161906 82102 162382 82170
rect 161906 82046 161930 82102
rect 161986 82046 162054 82102
rect 162110 82046 162178 82102
rect 162234 82046 162302 82102
rect 162358 82046 162382 82102
rect 161906 81978 162382 82046
rect 161906 81922 161930 81978
rect 161986 81922 162054 81978
rect 162110 81922 162178 81978
rect 162234 81922 162302 81978
rect 162358 81922 162382 81978
rect 161906 81888 162382 81922
rect 162738 82350 163358 99922
rect 162738 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 163358 82350
rect 162738 82226 163358 82294
rect 162738 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 163358 82226
rect 162738 82102 163358 82170
rect 162738 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 163358 82102
rect 162738 81978 163358 82046
rect 162738 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 163358 81978
rect 161106 76350 161582 76384
rect 161106 76294 161130 76350
rect 161186 76294 161254 76350
rect 161310 76294 161378 76350
rect 161434 76294 161502 76350
rect 161558 76294 161582 76350
rect 161106 76226 161582 76294
rect 161106 76170 161130 76226
rect 161186 76170 161254 76226
rect 161310 76170 161378 76226
rect 161434 76170 161502 76226
rect 161558 76170 161582 76226
rect 161106 76102 161582 76170
rect 161106 76046 161130 76102
rect 161186 76046 161254 76102
rect 161310 76046 161378 76102
rect 161434 76046 161502 76102
rect 161558 76046 161582 76102
rect 161106 75978 161582 76046
rect 161106 75922 161130 75978
rect 161186 75922 161254 75978
rect 161310 75922 161378 75978
rect 161434 75922 161502 75978
rect 161558 75922 161582 75978
rect 161106 75888 161582 75922
rect 161906 64350 162382 64384
rect 161906 64294 161930 64350
rect 161986 64294 162054 64350
rect 162110 64294 162178 64350
rect 162234 64294 162302 64350
rect 162358 64294 162382 64350
rect 161906 64226 162382 64294
rect 161906 64170 161930 64226
rect 161986 64170 162054 64226
rect 162110 64170 162178 64226
rect 162234 64170 162302 64226
rect 162358 64170 162382 64226
rect 161906 64102 162382 64170
rect 161906 64046 161930 64102
rect 161986 64046 162054 64102
rect 162110 64046 162178 64102
rect 162234 64046 162302 64102
rect 162358 64046 162382 64102
rect 161906 63978 162382 64046
rect 161906 63922 161930 63978
rect 161986 63922 162054 63978
rect 162110 63922 162178 63978
rect 162234 63922 162302 63978
rect 162358 63922 162382 63978
rect 161906 63888 162382 63922
rect 162738 64350 163358 81922
rect 162738 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 163358 64350
rect 162738 64226 163358 64294
rect 162738 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 163358 64226
rect 162738 64102 163358 64170
rect 162738 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 163358 64102
rect 162738 63978 163358 64046
rect 162738 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 163358 63978
rect 161106 58350 161582 58384
rect 161106 58294 161130 58350
rect 161186 58294 161254 58350
rect 161310 58294 161378 58350
rect 161434 58294 161502 58350
rect 161558 58294 161582 58350
rect 161106 58226 161582 58294
rect 161106 58170 161130 58226
rect 161186 58170 161254 58226
rect 161310 58170 161378 58226
rect 161434 58170 161502 58226
rect 161558 58170 161582 58226
rect 161106 58102 161582 58170
rect 161106 58046 161130 58102
rect 161186 58046 161254 58102
rect 161310 58046 161378 58102
rect 161434 58046 161502 58102
rect 161558 58046 161582 58102
rect 161106 57978 161582 58046
rect 161106 57922 161130 57978
rect 161186 57922 161254 57978
rect 161310 57922 161378 57978
rect 161434 57922 161502 57978
rect 161558 57922 161582 57978
rect 161106 57888 161582 57922
rect 161906 46350 162382 46384
rect 161906 46294 161930 46350
rect 161986 46294 162054 46350
rect 162110 46294 162178 46350
rect 162234 46294 162302 46350
rect 162358 46294 162382 46350
rect 161906 46226 162382 46294
rect 161906 46170 161930 46226
rect 161986 46170 162054 46226
rect 162110 46170 162178 46226
rect 162234 46170 162302 46226
rect 162358 46170 162382 46226
rect 161906 46102 162382 46170
rect 161906 46046 161930 46102
rect 161986 46046 162054 46102
rect 162110 46046 162178 46102
rect 162234 46046 162302 46102
rect 162358 46046 162382 46102
rect 161906 45978 162382 46046
rect 161906 45922 161930 45978
rect 161986 45922 162054 45978
rect 162110 45922 162178 45978
rect 162234 45922 162302 45978
rect 162358 45922 162382 45978
rect 161906 45888 162382 45922
rect 162738 46350 163358 63922
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 160412 4274 160468 4284
rect 162738 28350 163358 45922
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 162738 10350 163358 27922
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 143612 4050 143668 4060
rect 159018 4102 159638 4170
rect 137228 3378 137284 3388
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 -1120 163358 9922
rect 167916 4228 167972 170522
rect 168812 145684 168868 286524
rect 173068 285684 173124 285694
rect 168812 145618 168868 145628
rect 171276 281428 171332 281438
rect 167916 4162 167972 4172
rect 171276 4228 171332 281372
rect 171968 190350 172288 190384
rect 171968 190294 172038 190350
rect 172094 190294 172162 190350
rect 172218 190294 172288 190350
rect 171968 190226 172288 190294
rect 171968 190170 172038 190226
rect 172094 190170 172162 190226
rect 172218 190170 172288 190226
rect 171968 190102 172288 190170
rect 171968 190046 172038 190102
rect 172094 190046 172162 190102
rect 172218 190046 172288 190102
rect 171968 189978 172288 190046
rect 171968 189922 172038 189978
rect 172094 189922 172162 189978
rect 172218 189922 172288 189978
rect 171968 189888 172288 189922
rect 171968 172350 172288 172384
rect 171968 172294 172038 172350
rect 172094 172294 172162 172350
rect 172218 172294 172288 172350
rect 171968 172226 172288 172294
rect 171968 172170 172038 172226
rect 172094 172170 172162 172226
rect 172218 172170 172288 172226
rect 171968 172102 172288 172170
rect 171968 172046 172038 172102
rect 172094 172046 172162 172102
rect 172218 172046 172288 172102
rect 171968 171978 172288 172046
rect 171968 171922 172038 171978
rect 172094 171922 172162 171978
rect 172218 171922 172288 171978
rect 171968 171888 172288 171922
rect 173068 144004 173124 285628
rect 174748 285684 174804 285694
rect 174748 145796 174804 285628
rect 174748 145730 174804 145740
rect 173068 143938 173124 143948
rect 177212 143668 177268 286860
rect 178108 285684 178164 285694
rect 178108 143892 178164 285628
rect 178108 143826 178164 143836
rect 179676 158788 179732 158798
rect 177212 143602 177268 143612
rect 171276 4162 171332 4172
rect 179676 4116 179732 158732
rect 180572 148708 180628 286972
rect 183148 285684 183204 285694
rect 180572 148642 180628 148652
rect 182252 210868 182308 210878
rect 179676 4050 179732 4060
rect 180572 143668 180628 143678
rect 180572 3892 180628 143612
rect 182252 4116 182308 210812
rect 183148 143780 183204 285628
rect 184828 285684 184884 285694
rect 184828 157108 184884 285628
rect 188188 285684 188244 285694
rect 187328 202350 187648 202384
rect 187328 202294 187398 202350
rect 187454 202294 187522 202350
rect 187578 202294 187648 202350
rect 187328 202226 187648 202294
rect 187328 202170 187398 202226
rect 187454 202170 187522 202226
rect 187578 202170 187648 202226
rect 187328 202102 187648 202170
rect 187328 202046 187398 202102
rect 187454 202046 187522 202102
rect 187578 202046 187648 202102
rect 187328 201978 187648 202046
rect 187328 201922 187398 201978
rect 187454 201922 187522 201978
rect 187578 201922 187648 201978
rect 187328 201888 187648 201922
rect 187328 184350 187648 184384
rect 187328 184294 187398 184350
rect 187454 184294 187522 184350
rect 187578 184294 187648 184350
rect 187328 184226 187648 184294
rect 187328 184170 187398 184226
rect 187454 184170 187522 184226
rect 187578 184170 187648 184226
rect 187328 184102 187648 184170
rect 187328 184046 187398 184102
rect 187454 184046 187522 184102
rect 187578 184046 187648 184102
rect 187328 183978 187648 184046
rect 187328 183922 187398 183978
rect 187454 183922 187522 183978
rect 187578 183922 187648 183978
rect 187328 183888 187648 183922
rect 184828 157042 184884 157052
rect 185612 175618 185668 175628
rect 183148 143714 183204 143724
rect 185612 4228 185668 175562
rect 187328 166350 187648 166384
rect 187328 166294 187398 166350
rect 187454 166294 187522 166350
rect 187578 166294 187648 166350
rect 187328 166226 187648 166294
rect 187328 166170 187398 166226
rect 187454 166170 187522 166226
rect 187578 166170 187648 166226
rect 187328 166102 187648 166170
rect 187328 166046 187398 166102
rect 187454 166046 187522 166102
rect 187578 166046 187648 166102
rect 187328 165978 187648 166046
rect 187328 165922 187398 165978
rect 187454 165922 187522 165978
rect 187578 165922 187648 165978
rect 187328 165888 187648 165922
rect 188188 150612 188244 285628
rect 189738 274350 190358 291922
rect 193458 298350 194078 299890
rect 193458 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 194078 298350
rect 193458 298226 194078 298294
rect 193458 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 194078 298226
rect 193458 298102 194078 298170
rect 193458 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 194078 298102
rect 193458 297978 194078 298046
rect 193458 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 194078 297978
rect 189738 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 190358 274350
rect 189738 274226 190358 274294
rect 189738 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 190358 274226
rect 189738 274102 190358 274170
rect 189738 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 190358 274102
rect 189738 273978 190358 274046
rect 189738 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 190358 273978
rect 189738 256350 190358 273922
rect 189738 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 190358 256350
rect 189738 256226 190358 256294
rect 189738 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 190358 256226
rect 189738 256102 190358 256170
rect 189738 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 190358 256102
rect 189738 255978 190358 256046
rect 189738 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 190358 255978
rect 189738 238350 190358 255922
rect 189738 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 190358 238350
rect 189738 238226 190358 238294
rect 189738 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 190358 238226
rect 189738 238102 190358 238170
rect 189738 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 190358 238102
rect 189738 237978 190358 238046
rect 189738 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 190358 237978
rect 189738 220350 190358 237922
rect 189738 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 190358 220350
rect 189738 220226 190358 220294
rect 189738 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 190358 220226
rect 189738 220102 190358 220170
rect 189738 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 190358 220102
rect 189738 219978 190358 220046
rect 189738 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 190358 219978
rect 189738 202350 190358 219922
rect 189738 202294 189834 202350
rect 189890 202294 189958 202350
rect 190014 202294 190082 202350
rect 190138 202294 190206 202350
rect 190262 202294 190358 202350
rect 189738 202226 190358 202294
rect 189738 202170 189834 202226
rect 189890 202170 189958 202226
rect 190014 202170 190082 202226
rect 190138 202170 190206 202226
rect 190262 202170 190358 202226
rect 189738 202102 190358 202170
rect 189738 202046 189834 202102
rect 189890 202046 189958 202102
rect 190014 202046 190082 202102
rect 190138 202046 190206 202102
rect 190262 202046 190358 202102
rect 189738 201978 190358 202046
rect 189738 201922 189834 201978
rect 189890 201922 189958 201978
rect 190014 201922 190082 201978
rect 190138 201922 190206 201978
rect 190262 201922 190358 201978
rect 189738 184350 190358 201922
rect 189738 184294 189834 184350
rect 189890 184294 189958 184350
rect 190014 184294 190082 184350
rect 190138 184294 190206 184350
rect 190262 184294 190358 184350
rect 189738 184226 190358 184294
rect 189738 184170 189834 184226
rect 189890 184170 189958 184226
rect 190014 184170 190082 184226
rect 190138 184170 190206 184226
rect 190262 184170 190358 184226
rect 189738 184102 190358 184170
rect 189738 184046 189834 184102
rect 189890 184046 189958 184102
rect 190014 184046 190082 184102
rect 190138 184046 190206 184102
rect 190262 184046 190358 184102
rect 189738 183978 190358 184046
rect 189738 183922 189834 183978
rect 189890 183922 189958 183978
rect 190014 183922 190082 183978
rect 190138 183922 190206 183978
rect 190262 183922 190358 183978
rect 188188 150546 188244 150556
rect 188972 173998 189028 174008
rect 188972 4340 189028 173942
rect 188972 4274 189028 4284
rect 189738 166350 190358 183922
rect 189738 166294 189834 166350
rect 189890 166294 189958 166350
rect 190014 166294 190082 166350
rect 190138 166294 190206 166350
rect 190262 166294 190358 166350
rect 189738 166226 190358 166294
rect 189738 166170 189834 166226
rect 189890 166170 189958 166226
rect 190014 166170 190082 166226
rect 190138 166170 190206 166226
rect 190262 166170 190358 166226
rect 189738 166102 190358 166170
rect 189738 166046 189834 166102
rect 189890 166046 189958 166102
rect 190014 166046 190082 166102
rect 190138 166046 190206 166102
rect 190262 166046 190358 166102
rect 189738 165978 190358 166046
rect 189738 165922 189834 165978
rect 189890 165922 189958 165978
rect 190014 165922 190082 165978
rect 190138 165922 190206 165978
rect 190262 165922 190358 165978
rect 189738 148350 190358 165922
rect 191548 285684 191604 285694
rect 191548 158900 191604 285628
rect 193458 280350 194078 297922
rect 202688 298350 203008 298384
rect 202688 298294 202758 298350
rect 202814 298294 202882 298350
rect 202938 298294 203008 298350
rect 202688 298226 203008 298294
rect 202688 298170 202758 298226
rect 202814 298170 202882 298226
rect 202938 298170 203008 298226
rect 202688 298102 203008 298170
rect 202688 298046 202758 298102
rect 202814 298046 202882 298102
rect 202938 298046 203008 298102
rect 202688 297978 203008 298046
rect 202688 297922 202758 297978
rect 202814 297922 202882 297978
rect 202938 297922 203008 297978
rect 202688 297888 203008 297922
rect 220458 292350 221078 299890
rect 220458 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 221078 292350
rect 220458 292226 221078 292294
rect 220458 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 221078 292226
rect 220458 292102 221078 292170
rect 220458 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 221078 292102
rect 220458 291978 221078 292046
rect 220458 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 221078 291978
rect 200732 286468 200788 286478
rect 197372 285796 197428 285806
rect 193458 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 194078 280350
rect 193458 280226 194078 280294
rect 193458 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 194078 280226
rect 193458 280102 194078 280170
rect 193458 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 194078 280102
rect 193458 279978 194078 280046
rect 193458 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 194078 279978
rect 193458 262350 194078 279922
rect 193458 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 194078 262350
rect 193458 262226 194078 262294
rect 193458 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 194078 262226
rect 193458 262102 194078 262170
rect 193458 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 194078 262102
rect 193458 261978 194078 262046
rect 193458 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 194078 261978
rect 193458 244350 194078 261922
rect 193458 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 194078 244350
rect 193458 244226 194078 244294
rect 193458 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 194078 244226
rect 193458 244102 194078 244170
rect 193458 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 194078 244102
rect 193458 243978 194078 244046
rect 193458 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 194078 243978
rect 193458 226350 194078 243922
rect 193458 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 194078 226350
rect 193458 226226 194078 226294
rect 193458 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 194078 226226
rect 193458 226102 194078 226170
rect 193458 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 194078 226102
rect 193458 225978 194078 226046
rect 193458 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 194078 225978
rect 193458 208350 194078 225922
rect 193458 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 194078 208350
rect 193458 208226 194078 208294
rect 193458 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 194078 208226
rect 193458 208102 194078 208170
rect 193458 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 194078 208102
rect 193458 207978 194078 208046
rect 193458 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 194078 207978
rect 193458 190350 194078 207922
rect 193458 190294 193554 190350
rect 193610 190294 193678 190350
rect 193734 190294 193802 190350
rect 193858 190294 193926 190350
rect 193982 190294 194078 190350
rect 193458 190226 194078 190294
rect 193458 190170 193554 190226
rect 193610 190170 193678 190226
rect 193734 190170 193802 190226
rect 193858 190170 193926 190226
rect 193982 190170 194078 190226
rect 193458 190102 194078 190170
rect 193458 190046 193554 190102
rect 193610 190046 193678 190102
rect 193734 190046 193802 190102
rect 193858 190046 193926 190102
rect 193982 190046 194078 190102
rect 193458 189978 194078 190046
rect 193458 189922 193554 189978
rect 193610 189922 193678 189978
rect 193734 189922 193802 189978
rect 193858 189922 193926 189978
rect 193982 189922 194078 189978
rect 193458 172350 194078 189922
rect 193458 172294 193554 172350
rect 193610 172294 193678 172350
rect 193734 172294 193802 172350
rect 193858 172294 193926 172350
rect 193982 172294 194078 172350
rect 193458 172226 194078 172294
rect 193458 172170 193554 172226
rect 193610 172170 193678 172226
rect 193734 172170 193802 172226
rect 193858 172170 193926 172226
rect 193982 172170 194078 172226
rect 193458 172102 194078 172170
rect 193458 172046 193554 172102
rect 193610 172046 193678 172102
rect 193734 172046 193802 172102
rect 193858 172046 193926 172102
rect 193982 172046 194078 172102
rect 193458 171978 194078 172046
rect 193458 171922 193554 171978
rect 193610 171922 193678 171978
rect 193734 171922 193802 171978
rect 193858 171922 193926 171978
rect 193982 171922 194078 171978
rect 191548 158834 191604 158844
rect 192332 170758 192388 170768
rect 189738 148294 189834 148350
rect 189890 148294 189958 148350
rect 190014 148294 190082 148350
rect 190138 148294 190206 148350
rect 190262 148294 190358 148350
rect 189738 148226 190358 148294
rect 189738 148170 189834 148226
rect 189890 148170 189958 148226
rect 190014 148170 190082 148226
rect 190138 148170 190206 148226
rect 190262 148170 190358 148226
rect 189738 148102 190358 148170
rect 189738 148046 189834 148102
rect 189890 148046 189958 148102
rect 190014 148046 190082 148102
rect 190138 148046 190206 148102
rect 190262 148046 190358 148102
rect 189738 147978 190358 148046
rect 189738 147922 189834 147978
rect 189890 147922 189958 147978
rect 190014 147922 190082 147978
rect 190138 147922 190206 147978
rect 190262 147922 190358 147978
rect 189738 130350 190358 147922
rect 189738 130294 189834 130350
rect 189890 130294 189958 130350
rect 190014 130294 190082 130350
rect 190138 130294 190206 130350
rect 190262 130294 190358 130350
rect 189738 130226 190358 130294
rect 189738 130170 189834 130226
rect 189890 130170 189958 130226
rect 190014 130170 190082 130226
rect 190138 130170 190206 130226
rect 190262 130170 190358 130226
rect 189738 130102 190358 130170
rect 189738 130046 189834 130102
rect 189890 130046 189958 130102
rect 190014 130046 190082 130102
rect 190138 130046 190206 130102
rect 190262 130046 190358 130102
rect 189738 129978 190358 130046
rect 189738 129922 189834 129978
rect 189890 129922 189958 129978
rect 190014 129922 190082 129978
rect 190138 129922 190206 129978
rect 190262 129922 190358 129978
rect 189738 112350 190358 129922
rect 189738 112294 189834 112350
rect 189890 112294 189958 112350
rect 190014 112294 190082 112350
rect 190138 112294 190206 112350
rect 190262 112294 190358 112350
rect 189738 112226 190358 112294
rect 189738 112170 189834 112226
rect 189890 112170 189958 112226
rect 190014 112170 190082 112226
rect 190138 112170 190206 112226
rect 190262 112170 190358 112226
rect 189738 112102 190358 112170
rect 189738 112046 189834 112102
rect 189890 112046 189958 112102
rect 190014 112046 190082 112102
rect 190138 112046 190206 112102
rect 190262 112046 190358 112102
rect 189738 111978 190358 112046
rect 189738 111922 189834 111978
rect 189890 111922 189958 111978
rect 190014 111922 190082 111978
rect 190138 111922 190206 111978
rect 190262 111922 190358 111978
rect 189738 94350 190358 111922
rect 189738 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 190358 94350
rect 189738 94226 190358 94294
rect 189738 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 190358 94226
rect 189738 94102 190358 94170
rect 189738 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 190358 94102
rect 189738 93978 190358 94046
rect 189738 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 190358 93978
rect 189738 76350 190358 93922
rect 189738 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 190358 76350
rect 189738 76226 190358 76294
rect 189738 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 190358 76226
rect 189738 76102 190358 76170
rect 189738 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 190358 76102
rect 189738 75978 190358 76046
rect 189738 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 190358 75978
rect 189738 58350 190358 75922
rect 189738 58294 189834 58350
rect 189890 58294 189958 58350
rect 190014 58294 190082 58350
rect 190138 58294 190206 58350
rect 190262 58294 190358 58350
rect 189738 58226 190358 58294
rect 189738 58170 189834 58226
rect 189890 58170 189958 58226
rect 190014 58170 190082 58226
rect 190138 58170 190206 58226
rect 190262 58170 190358 58226
rect 189738 58102 190358 58170
rect 189738 58046 189834 58102
rect 189890 58046 189958 58102
rect 190014 58046 190082 58102
rect 190138 58046 190206 58102
rect 190262 58046 190358 58102
rect 189738 57978 190358 58046
rect 189738 57922 189834 57978
rect 189890 57922 189958 57978
rect 190014 57922 190082 57978
rect 190138 57922 190206 57978
rect 190262 57922 190358 57978
rect 189738 40350 190358 57922
rect 189738 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 190358 40350
rect 189738 40226 190358 40294
rect 189738 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 190358 40226
rect 189738 40102 190358 40170
rect 189738 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 190358 40102
rect 189738 39978 190358 40046
rect 189738 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 190358 39978
rect 189738 22350 190358 39922
rect 189738 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 190358 22350
rect 189738 22226 190358 22294
rect 189738 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 190358 22226
rect 189738 22102 190358 22170
rect 189738 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 190358 22102
rect 189738 21978 190358 22046
rect 189738 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 190358 21978
rect 189738 4350 190358 21922
rect 192332 4564 192388 170702
rect 192332 4498 192388 4508
rect 193458 154350 194078 171922
rect 193458 154294 193554 154350
rect 193610 154294 193678 154350
rect 193734 154294 193802 154350
rect 193858 154294 193926 154350
rect 193982 154294 194078 154350
rect 193458 154226 194078 154294
rect 193458 154170 193554 154226
rect 193610 154170 193678 154226
rect 193734 154170 193802 154226
rect 193858 154170 193926 154226
rect 193982 154170 194078 154226
rect 193458 154102 194078 154170
rect 193458 154046 193554 154102
rect 193610 154046 193678 154102
rect 193734 154046 193802 154102
rect 193858 154046 193926 154102
rect 193982 154046 194078 154102
rect 193458 153978 194078 154046
rect 193458 153922 193554 153978
rect 193610 153922 193678 153978
rect 193734 153922 193802 153978
rect 193858 153922 193926 153978
rect 193982 153922 194078 153978
rect 193458 136350 194078 153922
rect 194908 285684 194964 285694
rect 194908 145460 194964 285628
rect 194908 145394 194964 145404
rect 195692 168958 195748 168968
rect 193458 136294 193554 136350
rect 193610 136294 193678 136350
rect 193734 136294 193802 136350
rect 193858 136294 193926 136350
rect 193982 136294 194078 136350
rect 193458 136226 194078 136294
rect 193458 136170 193554 136226
rect 193610 136170 193678 136226
rect 193734 136170 193802 136226
rect 193858 136170 193926 136226
rect 193982 136170 194078 136226
rect 193458 136102 194078 136170
rect 193458 136046 193554 136102
rect 193610 136046 193678 136102
rect 193734 136046 193802 136102
rect 193858 136046 193926 136102
rect 193982 136046 194078 136102
rect 193458 135978 194078 136046
rect 193458 135922 193554 135978
rect 193610 135922 193678 135978
rect 193734 135922 193802 135978
rect 193858 135922 193926 135978
rect 193982 135922 194078 135978
rect 193458 118350 194078 135922
rect 193458 118294 193554 118350
rect 193610 118294 193678 118350
rect 193734 118294 193802 118350
rect 193858 118294 193926 118350
rect 193982 118294 194078 118350
rect 193458 118226 194078 118294
rect 193458 118170 193554 118226
rect 193610 118170 193678 118226
rect 193734 118170 193802 118226
rect 193858 118170 193926 118226
rect 193982 118170 194078 118226
rect 193458 118102 194078 118170
rect 193458 118046 193554 118102
rect 193610 118046 193678 118102
rect 193734 118046 193802 118102
rect 193858 118046 193926 118102
rect 193982 118046 194078 118102
rect 193458 117978 194078 118046
rect 193458 117922 193554 117978
rect 193610 117922 193678 117978
rect 193734 117922 193802 117978
rect 193858 117922 193926 117978
rect 193982 117922 194078 117978
rect 193458 100350 194078 117922
rect 193458 100294 193554 100350
rect 193610 100294 193678 100350
rect 193734 100294 193802 100350
rect 193858 100294 193926 100350
rect 193982 100294 194078 100350
rect 193458 100226 194078 100294
rect 193458 100170 193554 100226
rect 193610 100170 193678 100226
rect 193734 100170 193802 100226
rect 193858 100170 193926 100226
rect 193982 100170 194078 100226
rect 193458 100102 194078 100170
rect 193458 100046 193554 100102
rect 193610 100046 193678 100102
rect 193734 100046 193802 100102
rect 193858 100046 193926 100102
rect 193982 100046 194078 100102
rect 193458 99978 194078 100046
rect 193458 99922 193554 99978
rect 193610 99922 193678 99978
rect 193734 99922 193802 99978
rect 193858 99922 193926 99978
rect 193982 99922 194078 99978
rect 193458 82350 194078 99922
rect 193458 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 194078 82350
rect 193458 82226 194078 82294
rect 193458 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 194078 82226
rect 193458 82102 194078 82170
rect 193458 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 194078 82102
rect 193458 81978 194078 82046
rect 193458 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 194078 81978
rect 193458 64350 194078 81922
rect 193458 64294 193554 64350
rect 193610 64294 193678 64350
rect 193734 64294 193802 64350
rect 193858 64294 193926 64350
rect 193982 64294 194078 64350
rect 193458 64226 194078 64294
rect 193458 64170 193554 64226
rect 193610 64170 193678 64226
rect 193734 64170 193802 64226
rect 193858 64170 193926 64226
rect 193982 64170 194078 64226
rect 193458 64102 194078 64170
rect 193458 64046 193554 64102
rect 193610 64046 193678 64102
rect 193734 64046 193802 64102
rect 193858 64046 193926 64102
rect 193982 64046 194078 64102
rect 193458 63978 194078 64046
rect 193458 63922 193554 63978
rect 193610 63922 193678 63978
rect 193734 63922 193802 63978
rect 193858 63922 193926 63978
rect 193982 63922 194078 63978
rect 193458 46350 194078 63922
rect 193458 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 194078 46350
rect 193458 46226 194078 46294
rect 193458 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 194078 46226
rect 193458 46102 194078 46170
rect 193458 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 194078 46102
rect 193458 45978 194078 46046
rect 193458 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 194078 45978
rect 193458 28350 194078 45922
rect 193458 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 194078 28350
rect 193458 28226 194078 28294
rect 193458 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 194078 28226
rect 193458 28102 194078 28170
rect 193458 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 194078 28102
rect 193458 27978 194078 28046
rect 193458 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 194078 27978
rect 193458 10350 194078 27922
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 185612 4162 185668 4172
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 182252 4050 182308 4060
rect 189738 4102 190358 4170
rect 180572 3826 180628 3836
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 -1120 194078 9922
rect 195692 4452 195748 168902
rect 197372 147252 197428 285740
rect 198268 285684 198324 285694
rect 198268 167338 198324 285628
rect 200732 170578 200788 286412
rect 203308 285684 203364 285694
rect 202688 190350 203008 190384
rect 202688 190294 202758 190350
rect 202814 190294 202882 190350
rect 202938 190294 203008 190350
rect 202688 190226 203008 190294
rect 202688 190170 202758 190226
rect 202814 190170 202882 190226
rect 202938 190170 203008 190226
rect 202688 190102 203008 190170
rect 202688 190046 202758 190102
rect 202814 190046 202882 190102
rect 202938 190046 203008 190102
rect 202688 189978 203008 190046
rect 202688 189922 202758 189978
rect 202814 189922 202882 189978
rect 202938 189922 203008 189978
rect 202688 189888 203008 189922
rect 203308 173818 203364 285628
rect 203308 173752 203364 173762
rect 208348 285684 208404 285694
rect 202688 172350 203008 172384
rect 202688 172294 202758 172350
rect 202814 172294 202882 172350
rect 202938 172294 203008 172350
rect 202688 172226 203008 172294
rect 202688 172170 202758 172226
rect 202814 172170 202882 172226
rect 202938 172170 203008 172226
rect 202688 172102 203008 172170
rect 202688 172046 202758 172102
rect 202814 172046 202882 172102
rect 202938 172046 203008 172102
rect 202688 171978 203008 172046
rect 202688 171922 202758 171978
rect 202814 171922 202882 171978
rect 202938 171922 203008 171978
rect 202688 171888 203008 171922
rect 200732 170512 200788 170522
rect 208348 168778 208404 285628
rect 213388 285684 213444 285694
rect 213388 168958 213444 285628
rect 215068 285684 215124 285694
rect 215068 170758 215124 285628
rect 218428 285684 218484 285694
rect 218048 202350 218368 202384
rect 218048 202294 218118 202350
rect 218174 202294 218242 202350
rect 218298 202294 218368 202350
rect 218048 202226 218368 202294
rect 218048 202170 218118 202226
rect 218174 202170 218242 202226
rect 218298 202170 218368 202226
rect 218048 202102 218368 202170
rect 218048 202046 218118 202102
rect 218174 202046 218242 202102
rect 218298 202046 218368 202102
rect 218048 201978 218368 202046
rect 218048 201922 218118 201978
rect 218174 201922 218242 201978
rect 218298 201922 218368 201978
rect 218048 201888 218368 201922
rect 218048 184350 218368 184384
rect 218048 184294 218118 184350
rect 218174 184294 218242 184350
rect 218298 184294 218368 184350
rect 218048 184226 218368 184294
rect 218048 184170 218118 184226
rect 218174 184170 218242 184226
rect 218298 184170 218368 184226
rect 218048 184102 218368 184170
rect 218048 184046 218118 184102
rect 218174 184046 218242 184102
rect 218298 184046 218368 184102
rect 218048 183978 218368 184046
rect 218048 183922 218118 183978
rect 218174 183922 218242 183978
rect 218298 183922 218368 183978
rect 218048 183888 218368 183922
rect 218428 175618 218484 285628
rect 218428 175552 218484 175562
rect 220458 274350 221078 291922
rect 224178 298350 224798 299890
rect 224178 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 224798 298350
rect 224178 298226 224798 298294
rect 224178 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 224798 298226
rect 224178 298102 224798 298170
rect 224178 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 224798 298102
rect 224178 297978 224798 298046
rect 224178 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 224798 297978
rect 220458 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 221078 274350
rect 220458 274226 221078 274294
rect 220458 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 221078 274226
rect 220458 274102 221078 274170
rect 220458 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 221078 274102
rect 220458 273978 221078 274046
rect 220458 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 221078 273978
rect 220458 256350 221078 273922
rect 220458 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 221078 256350
rect 220458 256226 221078 256294
rect 220458 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 221078 256226
rect 220458 256102 221078 256170
rect 220458 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 221078 256102
rect 220458 255978 221078 256046
rect 220458 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 221078 255978
rect 220458 238350 221078 255922
rect 220458 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 221078 238350
rect 220458 238226 221078 238294
rect 220458 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 221078 238226
rect 220458 238102 221078 238170
rect 220458 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 221078 238102
rect 220458 237978 221078 238046
rect 220458 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 221078 237978
rect 220458 220350 221078 237922
rect 220458 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 221078 220350
rect 220458 220226 221078 220294
rect 220458 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 221078 220226
rect 220458 220102 221078 220170
rect 220458 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 221078 220102
rect 220458 219978 221078 220046
rect 220458 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 221078 219978
rect 220458 202350 221078 219922
rect 220458 202294 220554 202350
rect 220610 202294 220678 202350
rect 220734 202294 220802 202350
rect 220858 202294 220926 202350
rect 220982 202294 221078 202350
rect 220458 202226 221078 202294
rect 220458 202170 220554 202226
rect 220610 202170 220678 202226
rect 220734 202170 220802 202226
rect 220858 202170 220926 202226
rect 220982 202170 221078 202226
rect 220458 202102 221078 202170
rect 220458 202046 220554 202102
rect 220610 202046 220678 202102
rect 220734 202046 220802 202102
rect 220858 202046 220926 202102
rect 220982 202046 221078 202102
rect 220458 201978 221078 202046
rect 220458 201922 220554 201978
rect 220610 201922 220678 201978
rect 220734 201922 220802 201978
rect 220858 201922 220926 201978
rect 220982 201922 221078 201978
rect 220458 184350 221078 201922
rect 220458 184294 220554 184350
rect 220610 184294 220678 184350
rect 220734 184294 220802 184350
rect 220858 184294 220926 184350
rect 220982 184294 221078 184350
rect 220458 184226 221078 184294
rect 220458 184170 220554 184226
rect 220610 184170 220678 184226
rect 220734 184170 220802 184226
rect 220858 184170 220926 184226
rect 220982 184170 221078 184226
rect 220458 184102 221078 184170
rect 220458 184046 220554 184102
rect 220610 184046 220678 184102
rect 220734 184046 220802 184102
rect 220858 184046 220926 184102
rect 220982 184046 221078 184102
rect 220458 183978 221078 184046
rect 220458 183922 220554 183978
rect 220610 183922 220678 183978
rect 220734 183922 220802 183978
rect 220858 183922 220926 183978
rect 220982 183922 221078 183978
rect 215068 170692 215124 170702
rect 220458 169150 221078 183922
rect 221788 285684 221844 285694
rect 221788 173998 221844 285628
rect 221788 173932 221844 173942
rect 224178 280350 224798 297922
rect 233408 298350 233728 298384
rect 233408 298294 233478 298350
rect 233534 298294 233602 298350
rect 233658 298294 233728 298350
rect 233408 298226 233728 298294
rect 233408 298170 233478 298226
rect 233534 298170 233602 298226
rect 233658 298170 233728 298226
rect 233408 298102 233728 298170
rect 233408 298046 233478 298102
rect 233534 298046 233602 298102
rect 233658 298046 233728 298102
rect 233408 297978 233728 298046
rect 233408 297922 233478 297978
rect 233534 297922 233602 297978
rect 233658 297922 233728 297978
rect 233408 297888 233728 297922
rect 251178 292350 251798 299890
rect 251178 292294 251274 292350
rect 251330 292294 251398 292350
rect 251454 292294 251522 292350
rect 251578 292294 251646 292350
rect 251702 292294 251798 292350
rect 251178 292226 251798 292294
rect 251178 292170 251274 292226
rect 251330 292170 251398 292226
rect 251454 292170 251522 292226
rect 251578 292170 251646 292226
rect 251702 292170 251798 292226
rect 251178 292102 251798 292170
rect 251178 292046 251274 292102
rect 251330 292046 251398 292102
rect 251454 292046 251522 292102
rect 251578 292046 251646 292102
rect 251702 292046 251798 292102
rect 251178 291978 251798 292046
rect 251178 291922 251274 291978
rect 251330 291922 251398 291978
rect 251454 291922 251522 291978
rect 251578 291922 251646 291978
rect 251702 291922 251798 291978
rect 247772 291508 247828 291518
rect 245196 289828 245252 289838
rect 230972 286468 231028 286478
rect 227612 285796 227668 285806
rect 224178 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 224798 280350
rect 224178 280226 224798 280294
rect 224178 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 224798 280226
rect 224178 280102 224798 280170
rect 224178 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 224798 280102
rect 224178 279978 224798 280046
rect 224178 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 224798 279978
rect 224178 262350 224798 279922
rect 224178 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 224798 262350
rect 224178 262226 224798 262294
rect 224178 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 224798 262226
rect 224178 262102 224798 262170
rect 224178 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 224798 262102
rect 224178 261978 224798 262046
rect 224178 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 224798 261978
rect 224178 244350 224798 261922
rect 224178 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 224798 244350
rect 224178 244226 224798 244294
rect 224178 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 224798 244226
rect 224178 244102 224798 244170
rect 224178 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 224798 244102
rect 224178 243978 224798 244046
rect 224178 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 224798 243978
rect 224178 226350 224798 243922
rect 224178 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 224798 226350
rect 224178 226226 224798 226294
rect 224178 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 224798 226226
rect 224178 226102 224798 226170
rect 224178 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 224798 226102
rect 224178 225978 224798 226046
rect 224178 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 224798 225978
rect 224178 208350 224798 225922
rect 224178 208294 224274 208350
rect 224330 208294 224398 208350
rect 224454 208294 224522 208350
rect 224578 208294 224646 208350
rect 224702 208294 224798 208350
rect 224178 208226 224798 208294
rect 224178 208170 224274 208226
rect 224330 208170 224398 208226
rect 224454 208170 224522 208226
rect 224578 208170 224646 208226
rect 224702 208170 224798 208226
rect 224178 208102 224798 208170
rect 224178 208046 224274 208102
rect 224330 208046 224398 208102
rect 224454 208046 224522 208102
rect 224578 208046 224646 208102
rect 224702 208046 224798 208102
rect 224178 207978 224798 208046
rect 224178 207922 224274 207978
rect 224330 207922 224398 207978
rect 224454 207922 224522 207978
rect 224578 207922 224646 207978
rect 224702 207922 224798 207978
rect 224178 190350 224798 207922
rect 224178 190294 224274 190350
rect 224330 190294 224398 190350
rect 224454 190294 224522 190350
rect 224578 190294 224646 190350
rect 224702 190294 224798 190350
rect 224178 190226 224798 190294
rect 224178 190170 224274 190226
rect 224330 190170 224398 190226
rect 224454 190170 224522 190226
rect 224578 190170 224646 190226
rect 224702 190170 224798 190226
rect 224178 190102 224798 190170
rect 224178 190046 224274 190102
rect 224330 190046 224398 190102
rect 224454 190046 224522 190102
rect 224578 190046 224646 190102
rect 224702 190046 224798 190102
rect 224178 189978 224798 190046
rect 224178 189922 224274 189978
rect 224330 189922 224398 189978
rect 224454 189922 224522 189978
rect 224578 189922 224646 189978
rect 224702 189922 224798 189978
rect 224178 172350 224798 189922
rect 224178 172294 224274 172350
rect 224330 172294 224398 172350
rect 224454 172294 224522 172350
rect 224578 172294 224646 172350
rect 224702 172294 224798 172350
rect 224178 172226 224798 172294
rect 224178 172170 224274 172226
rect 224330 172170 224398 172226
rect 224454 172170 224522 172226
rect 224578 172170 224646 172226
rect 224702 172170 224798 172226
rect 224178 172102 224798 172170
rect 224178 172046 224274 172102
rect 224330 172046 224398 172102
rect 224454 172046 224522 172102
rect 224578 172046 224646 172102
rect 224702 172046 224798 172102
rect 224178 171978 224798 172046
rect 224178 171922 224274 171978
rect 224330 171922 224398 171978
rect 224454 171922 224522 171978
rect 224578 171922 224646 171978
rect 224702 171922 224798 171978
rect 224178 169150 224798 171922
rect 225148 285684 225204 285694
rect 213388 168892 213444 168902
rect 208348 168712 208404 168722
rect 198268 167272 198324 167282
rect 218048 166350 218368 166384
rect 218048 166294 218118 166350
rect 218174 166294 218242 166350
rect 218298 166294 218368 166350
rect 218048 166226 218368 166294
rect 218048 166170 218118 166226
rect 218174 166170 218242 166226
rect 218298 166170 218368 166226
rect 218048 166102 218368 166170
rect 218048 166046 218118 166102
rect 218174 166046 218242 166102
rect 218298 166046 218368 166102
rect 218048 165978 218368 166046
rect 218048 165922 218118 165978
rect 218174 165922 218242 165978
rect 218298 165922 218368 165978
rect 218048 165888 218368 165922
rect 197372 147186 197428 147196
rect 220458 148350 221078 162274
rect 220458 148294 220554 148350
rect 220610 148294 220678 148350
rect 220734 148294 220802 148350
rect 220858 148294 220926 148350
rect 220982 148294 221078 148350
rect 220458 148226 221078 148294
rect 220458 148170 220554 148226
rect 220610 148170 220678 148226
rect 220734 148170 220802 148226
rect 220858 148170 220926 148226
rect 220982 148170 221078 148226
rect 220458 148102 221078 148170
rect 220458 148046 220554 148102
rect 220610 148046 220678 148102
rect 220734 148046 220802 148102
rect 220858 148046 220926 148102
rect 220982 148046 221078 148102
rect 220458 147978 221078 148046
rect 220458 147922 220554 147978
rect 220610 147922 220678 147978
rect 220734 147922 220802 147978
rect 220858 147922 220926 147978
rect 220982 147922 221078 147978
rect 219324 141958 219380 141968
rect 214620 141204 214676 141214
rect 214620 141058 214676 141148
rect 219324 141204 219380 141902
rect 219324 141138 219380 141148
rect 214620 140992 214676 141002
rect 195692 4386 195748 4396
rect 220458 130350 221078 147922
rect 220458 130294 220554 130350
rect 220610 130294 220678 130350
rect 220734 130294 220802 130350
rect 220858 130294 220926 130350
rect 220982 130294 221078 130350
rect 220458 130226 221078 130294
rect 220458 130170 220554 130226
rect 220610 130170 220678 130226
rect 220734 130170 220802 130226
rect 220858 130170 220926 130226
rect 220982 130170 221078 130226
rect 220458 130102 221078 130170
rect 220458 130046 220554 130102
rect 220610 130046 220678 130102
rect 220734 130046 220802 130102
rect 220858 130046 220926 130102
rect 220982 130046 221078 130102
rect 220458 129978 221078 130046
rect 220458 129922 220554 129978
rect 220610 129922 220678 129978
rect 220734 129922 220802 129978
rect 220858 129922 220926 129978
rect 220982 129922 221078 129978
rect 220458 112350 221078 129922
rect 220458 112294 220554 112350
rect 220610 112294 220678 112350
rect 220734 112294 220802 112350
rect 220858 112294 220926 112350
rect 220982 112294 221078 112350
rect 220458 112226 221078 112294
rect 220458 112170 220554 112226
rect 220610 112170 220678 112226
rect 220734 112170 220802 112226
rect 220858 112170 220926 112226
rect 220982 112170 221078 112226
rect 220458 112102 221078 112170
rect 220458 112046 220554 112102
rect 220610 112046 220678 112102
rect 220734 112046 220802 112102
rect 220858 112046 220926 112102
rect 220982 112046 221078 112102
rect 220458 111978 221078 112046
rect 220458 111922 220554 111978
rect 220610 111922 220678 111978
rect 220734 111922 220802 111978
rect 220858 111922 220926 111978
rect 220982 111922 221078 111978
rect 220458 94350 221078 111922
rect 220458 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 221078 94350
rect 220458 94226 221078 94294
rect 220458 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 221078 94226
rect 220458 94102 221078 94170
rect 220458 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 221078 94102
rect 220458 93978 221078 94046
rect 220458 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 221078 93978
rect 220458 76350 221078 93922
rect 220458 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 221078 76350
rect 220458 76226 221078 76294
rect 220458 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 221078 76226
rect 220458 76102 221078 76170
rect 220458 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 221078 76102
rect 220458 75978 221078 76046
rect 220458 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 221078 75978
rect 220458 58350 221078 75922
rect 220458 58294 220554 58350
rect 220610 58294 220678 58350
rect 220734 58294 220802 58350
rect 220858 58294 220926 58350
rect 220982 58294 221078 58350
rect 220458 58226 221078 58294
rect 220458 58170 220554 58226
rect 220610 58170 220678 58226
rect 220734 58170 220802 58226
rect 220858 58170 220926 58226
rect 220982 58170 221078 58226
rect 220458 58102 221078 58170
rect 220458 58046 220554 58102
rect 220610 58046 220678 58102
rect 220734 58046 220802 58102
rect 220858 58046 220926 58102
rect 220982 58046 221078 58102
rect 220458 57978 221078 58046
rect 220458 57922 220554 57978
rect 220610 57922 220678 57978
rect 220734 57922 220802 57978
rect 220858 57922 220926 57978
rect 220982 57922 221078 57978
rect 220458 40350 221078 57922
rect 220458 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 221078 40350
rect 220458 40226 221078 40294
rect 220458 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 221078 40226
rect 220458 40102 221078 40170
rect 220458 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 221078 40102
rect 220458 39978 221078 40046
rect 220458 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 221078 39978
rect 220458 22350 221078 39922
rect 220458 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 221078 22350
rect 220458 22226 221078 22294
rect 220458 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 221078 22226
rect 220458 22102 221078 22170
rect 220458 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 221078 22102
rect 220458 21978 221078 22046
rect 220458 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 221078 21978
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 4350 221078 21922
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 154350 224798 162274
rect 224178 154294 224274 154350
rect 224330 154294 224398 154350
rect 224454 154294 224522 154350
rect 224578 154294 224646 154350
rect 224702 154294 224798 154350
rect 224178 154226 224798 154294
rect 224178 154170 224274 154226
rect 224330 154170 224398 154226
rect 224454 154170 224522 154226
rect 224578 154170 224646 154226
rect 224702 154170 224798 154226
rect 224178 154102 224798 154170
rect 224178 154046 224274 154102
rect 224330 154046 224398 154102
rect 224454 154046 224522 154102
rect 224578 154046 224646 154102
rect 224702 154046 224798 154102
rect 224178 153978 224798 154046
rect 224178 153922 224274 153978
rect 224330 153922 224398 153978
rect 224454 153922 224522 153978
rect 224578 153922 224646 153978
rect 224702 153922 224798 153978
rect 224178 136350 224798 153922
rect 225148 143668 225204 285628
rect 225148 143602 225204 143612
rect 226716 159012 226772 159022
rect 224178 136294 224274 136350
rect 224330 136294 224398 136350
rect 224454 136294 224522 136350
rect 224578 136294 224646 136350
rect 224702 136294 224798 136350
rect 224178 136226 224798 136294
rect 224178 136170 224274 136226
rect 224330 136170 224398 136226
rect 224454 136170 224522 136226
rect 224578 136170 224646 136226
rect 224702 136170 224798 136226
rect 224178 136102 224798 136170
rect 224178 136046 224274 136102
rect 224330 136046 224398 136102
rect 224454 136046 224522 136102
rect 224578 136046 224646 136102
rect 224702 136046 224798 136102
rect 224178 135978 224798 136046
rect 224178 135922 224274 135978
rect 224330 135922 224398 135978
rect 224454 135922 224522 135978
rect 224578 135922 224646 135978
rect 224702 135922 224798 135978
rect 224178 118350 224798 135922
rect 224178 118294 224274 118350
rect 224330 118294 224398 118350
rect 224454 118294 224522 118350
rect 224578 118294 224646 118350
rect 224702 118294 224798 118350
rect 224178 118226 224798 118294
rect 224178 118170 224274 118226
rect 224330 118170 224398 118226
rect 224454 118170 224522 118226
rect 224578 118170 224646 118226
rect 224702 118170 224798 118226
rect 224178 118102 224798 118170
rect 224178 118046 224274 118102
rect 224330 118046 224398 118102
rect 224454 118046 224522 118102
rect 224578 118046 224646 118102
rect 224702 118046 224798 118102
rect 224178 117978 224798 118046
rect 224178 117922 224274 117978
rect 224330 117922 224398 117978
rect 224454 117922 224522 117978
rect 224578 117922 224646 117978
rect 224702 117922 224798 117978
rect 224178 100350 224798 117922
rect 224178 100294 224274 100350
rect 224330 100294 224398 100350
rect 224454 100294 224522 100350
rect 224578 100294 224646 100350
rect 224702 100294 224798 100350
rect 224178 100226 224798 100294
rect 224178 100170 224274 100226
rect 224330 100170 224398 100226
rect 224454 100170 224522 100226
rect 224578 100170 224646 100226
rect 224702 100170 224798 100226
rect 224178 100102 224798 100170
rect 224178 100046 224274 100102
rect 224330 100046 224398 100102
rect 224454 100046 224522 100102
rect 224578 100046 224646 100102
rect 224702 100046 224798 100102
rect 224178 99978 224798 100046
rect 224178 99922 224274 99978
rect 224330 99922 224398 99978
rect 224454 99922 224522 99978
rect 224578 99922 224646 99978
rect 224702 99922 224798 99978
rect 224178 82350 224798 99922
rect 224178 82294 224274 82350
rect 224330 82294 224398 82350
rect 224454 82294 224522 82350
rect 224578 82294 224646 82350
rect 224702 82294 224798 82350
rect 224178 82226 224798 82294
rect 224178 82170 224274 82226
rect 224330 82170 224398 82226
rect 224454 82170 224522 82226
rect 224578 82170 224646 82226
rect 224702 82170 224798 82226
rect 224178 82102 224798 82170
rect 224178 82046 224274 82102
rect 224330 82046 224398 82102
rect 224454 82046 224522 82102
rect 224578 82046 224646 82102
rect 224702 82046 224798 82102
rect 224178 81978 224798 82046
rect 224178 81922 224274 81978
rect 224330 81922 224398 81978
rect 224454 81922 224522 81978
rect 224578 81922 224646 81978
rect 224702 81922 224798 81978
rect 224178 64350 224798 81922
rect 224178 64294 224274 64350
rect 224330 64294 224398 64350
rect 224454 64294 224522 64350
rect 224578 64294 224646 64350
rect 224702 64294 224798 64350
rect 224178 64226 224798 64294
rect 224178 64170 224274 64226
rect 224330 64170 224398 64226
rect 224454 64170 224522 64226
rect 224578 64170 224646 64226
rect 224702 64170 224798 64226
rect 224178 64102 224798 64170
rect 224178 64046 224274 64102
rect 224330 64046 224398 64102
rect 224454 64046 224522 64102
rect 224578 64046 224646 64102
rect 224702 64046 224798 64102
rect 224178 63978 224798 64046
rect 224178 63922 224274 63978
rect 224330 63922 224398 63978
rect 224454 63922 224522 63978
rect 224578 63922 224646 63978
rect 224702 63922 224798 63978
rect 224178 46350 224798 63922
rect 224178 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 224798 46350
rect 224178 46226 224798 46294
rect 224178 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 224798 46226
rect 224178 46102 224798 46170
rect 224178 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 224798 46102
rect 224178 45978 224798 46046
rect 224178 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 224798 45978
rect 224178 28350 224798 45922
rect 224178 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 224798 28350
rect 224178 28226 224798 28294
rect 224178 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 224798 28226
rect 224178 28102 224798 28170
rect 224178 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 224798 28102
rect 224178 27978 224798 28046
rect 224178 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 224798 27978
rect 224178 10350 224798 27922
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 224178 -1120 224798 9922
rect 226716 4116 226772 158956
rect 227612 14308 227668 285740
rect 228508 285684 228564 285694
rect 228508 152404 228564 285628
rect 228508 152338 228564 152348
rect 227612 14242 227668 14252
rect 230972 6132 231028 286412
rect 231868 285684 231924 285694
rect 231868 158788 231924 285628
rect 237692 285684 237748 285694
rect 233408 190350 233728 190384
rect 233408 190294 233478 190350
rect 233534 190294 233602 190350
rect 233658 190294 233728 190350
rect 233408 190226 233728 190294
rect 233408 190170 233478 190226
rect 233534 190170 233602 190226
rect 233658 190170 233728 190226
rect 233408 190102 233728 190170
rect 233408 190046 233478 190102
rect 233534 190046 233602 190102
rect 233658 190046 233728 190102
rect 233408 189978 233728 190046
rect 233408 189922 233478 189978
rect 233534 189922 233602 189978
rect 233658 189922 233728 189978
rect 233408 189888 233728 189922
rect 233408 172350 233728 172384
rect 233408 172294 233478 172350
rect 233534 172294 233602 172350
rect 233658 172294 233728 172350
rect 233408 172226 233728 172294
rect 233408 172170 233478 172226
rect 233534 172170 233602 172226
rect 233658 172170 233728 172226
rect 233408 172102 233728 172170
rect 233408 172046 233478 172102
rect 233534 172046 233602 172102
rect 233658 172046 233728 172102
rect 233408 171978 233728 172046
rect 233408 171922 233478 171978
rect 233534 171922 233602 171978
rect 233658 171922 233728 171978
rect 233408 171888 233728 171922
rect 231868 158722 231924 158732
rect 233436 160356 233492 160366
rect 230972 6066 231028 6076
rect 226716 4050 226772 4060
rect 233436 4116 233492 160300
rect 237692 12628 237748 285628
rect 237692 12562 237748 12572
rect 239372 285684 239428 285694
rect 239372 7700 239428 285628
rect 243516 285684 243572 285694
rect 243516 143892 243572 285628
rect 243516 143826 243572 143836
rect 244636 142138 244692 142148
rect 244636 141204 244692 142082
rect 244636 141138 244692 141148
rect 239372 7634 239428 7644
rect 245196 4228 245252 289772
rect 246876 285684 246932 285694
rect 246876 146244 246932 285628
rect 246876 146178 246932 146188
rect 245420 140878 245476 140888
rect 245420 140644 245476 140822
rect 245420 140578 245476 140588
rect 245788 130350 246264 130384
rect 245788 130294 245812 130350
rect 245868 130294 245936 130350
rect 245992 130294 246060 130350
rect 246116 130294 246184 130350
rect 246240 130294 246264 130350
rect 245788 130226 246264 130294
rect 245788 130170 245812 130226
rect 245868 130170 245936 130226
rect 245992 130170 246060 130226
rect 246116 130170 246184 130226
rect 246240 130170 246264 130226
rect 245788 130102 246264 130170
rect 245788 130046 245812 130102
rect 245868 130046 245936 130102
rect 245992 130046 246060 130102
rect 246116 130046 246184 130102
rect 246240 130046 246264 130102
rect 245788 129978 246264 130046
rect 245788 129922 245812 129978
rect 245868 129922 245936 129978
rect 245992 129922 246060 129978
rect 246116 129922 246184 129978
rect 246240 129922 246264 129978
rect 245788 129888 246264 129922
rect 246588 118350 247064 118384
rect 246588 118294 246612 118350
rect 246668 118294 246736 118350
rect 246792 118294 246860 118350
rect 246916 118294 246984 118350
rect 247040 118294 247064 118350
rect 246588 118226 247064 118294
rect 246588 118170 246612 118226
rect 246668 118170 246736 118226
rect 246792 118170 246860 118226
rect 246916 118170 246984 118226
rect 247040 118170 247064 118226
rect 246588 118102 247064 118170
rect 246588 118046 246612 118102
rect 246668 118046 246736 118102
rect 246792 118046 246860 118102
rect 246916 118046 246984 118102
rect 247040 118046 247064 118102
rect 246588 117978 247064 118046
rect 246588 117922 246612 117978
rect 246668 117922 246736 117978
rect 246792 117922 246860 117978
rect 246916 117922 246984 117978
rect 247040 117922 247064 117978
rect 246588 117888 247064 117922
rect 245788 112350 246264 112384
rect 245788 112294 245812 112350
rect 245868 112294 245936 112350
rect 245992 112294 246060 112350
rect 246116 112294 246184 112350
rect 246240 112294 246264 112350
rect 245788 112226 246264 112294
rect 245788 112170 245812 112226
rect 245868 112170 245936 112226
rect 245992 112170 246060 112226
rect 246116 112170 246184 112226
rect 246240 112170 246264 112226
rect 245788 112102 246264 112170
rect 245788 112046 245812 112102
rect 245868 112046 245936 112102
rect 245992 112046 246060 112102
rect 246116 112046 246184 112102
rect 246240 112046 246264 112102
rect 245788 111978 246264 112046
rect 245788 111922 245812 111978
rect 245868 111922 245936 111978
rect 245992 111922 246060 111978
rect 246116 111922 246184 111978
rect 246240 111922 246264 111978
rect 245788 111888 246264 111922
rect 246588 100350 247064 100384
rect 246588 100294 246612 100350
rect 246668 100294 246736 100350
rect 246792 100294 246860 100350
rect 246916 100294 246984 100350
rect 247040 100294 247064 100350
rect 246588 100226 247064 100294
rect 246588 100170 246612 100226
rect 246668 100170 246736 100226
rect 246792 100170 246860 100226
rect 246916 100170 246984 100226
rect 247040 100170 247064 100226
rect 246588 100102 247064 100170
rect 246588 100046 246612 100102
rect 246668 100046 246736 100102
rect 246792 100046 246860 100102
rect 246916 100046 246984 100102
rect 247040 100046 247064 100102
rect 246588 99978 247064 100046
rect 246588 99922 246612 99978
rect 246668 99922 246736 99978
rect 246792 99922 246860 99978
rect 246916 99922 246984 99978
rect 247040 99922 247064 99978
rect 246588 99888 247064 99922
rect 245788 94350 246264 94384
rect 245788 94294 245812 94350
rect 245868 94294 245936 94350
rect 245992 94294 246060 94350
rect 246116 94294 246184 94350
rect 246240 94294 246264 94350
rect 245788 94226 246264 94294
rect 245788 94170 245812 94226
rect 245868 94170 245936 94226
rect 245992 94170 246060 94226
rect 246116 94170 246184 94226
rect 246240 94170 246264 94226
rect 245788 94102 246264 94170
rect 245788 94046 245812 94102
rect 245868 94046 245936 94102
rect 245992 94046 246060 94102
rect 246116 94046 246184 94102
rect 246240 94046 246264 94102
rect 245788 93978 246264 94046
rect 245788 93922 245812 93978
rect 245868 93922 245936 93978
rect 245992 93922 246060 93978
rect 246116 93922 246184 93978
rect 246240 93922 246264 93978
rect 245788 93888 246264 93922
rect 246588 82350 247064 82384
rect 246588 82294 246612 82350
rect 246668 82294 246736 82350
rect 246792 82294 246860 82350
rect 246916 82294 246984 82350
rect 247040 82294 247064 82350
rect 246588 82226 247064 82294
rect 246588 82170 246612 82226
rect 246668 82170 246736 82226
rect 246792 82170 246860 82226
rect 246916 82170 246984 82226
rect 247040 82170 247064 82226
rect 246588 82102 247064 82170
rect 246588 82046 246612 82102
rect 246668 82046 246736 82102
rect 246792 82046 246860 82102
rect 246916 82046 246984 82102
rect 247040 82046 247064 82102
rect 246588 81978 247064 82046
rect 246588 81922 246612 81978
rect 246668 81922 246736 81978
rect 246792 81922 246860 81978
rect 246916 81922 246984 81978
rect 247040 81922 247064 81978
rect 246588 81888 247064 81922
rect 245788 76350 246264 76384
rect 245788 76294 245812 76350
rect 245868 76294 245936 76350
rect 245992 76294 246060 76350
rect 246116 76294 246184 76350
rect 246240 76294 246264 76350
rect 245788 76226 246264 76294
rect 245788 76170 245812 76226
rect 245868 76170 245936 76226
rect 245992 76170 246060 76226
rect 246116 76170 246184 76226
rect 246240 76170 246264 76226
rect 245788 76102 246264 76170
rect 245788 76046 245812 76102
rect 245868 76046 245936 76102
rect 245992 76046 246060 76102
rect 246116 76046 246184 76102
rect 246240 76046 246264 76102
rect 245788 75978 246264 76046
rect 245788 75922 245812 75978
rect 245868 75922 245936 75978
rect 245992 75922 246060 75978
rect 246116 75922 246184 75978
rect 246240 75922 246264 75978
rect 245788 75888 246264 75922
rect 246588 64350 247064 64384
rect 246588 64294 246612 64350
rect 246668 64294 246736 64350
rect 246792 64294 246860 64350
rect 246916 64294 246984 64350
rect 247040 64294 247064 64350
rect 246588 64226 247064 64294
rect 246588 64170 246612 64226
rect 246668 64170 246736 64226
rect 246792 64170 246860 64226
rect 246916 64170 246984 64226
rect 247040 64170 247064 64226
rect 246588 64102 247064 64170
rect 246588 64046 246612 64102
rect 246668 64046 246736 64102
rect 246792 64046 246860 64102
rect 246916 64046 246984 64102
rect 247040 64046 247064 64102
rect 246588 63978 247064 64046
rect 246588 63922 246612 63978
rect 246668 63922 246736 63978
rect 246792 63922 246860 63978
rect 246916 63922 246984 63978
rect 247040 63922 247064 63978
rect 246588 63888 247064 63922
rect 245788 58350 246264 58384
rect 245788 58294 245812 58350
rect 245868 58294 245936 58350
rect 245992 58294 246060 58350
rect 246116 58294 246184 58350
rect 246240 58294 246264 58350
rect 245788 58226 246264 58294
rect 245788 58170 245812 58226
rect 245868 58170 245936 58226
rect 245992 58170 246060 58226
rect 246116 58170 246184 58226
rect 246240 58170 246264 58226
rect 245788 58102 246264 58170
rect 245788 58046 245812 58102
rect 245868 58046 245936 58102
rect 245992 58046 246060 58102
rect 246116 58046 246184 58102
rect 246240 58046 246264 58102
rect 245788 57978 246264 58046
rect 245788 57922 245812 57978
rect 245868 57922 245936 57978
rect 245992 57922 246060 57978
rect 246116 57922 246184 57978
rect 246240 57922 246264 57978
rect 245788 57888 246264 57922
rect 246588 46350 247064 46384
rect 246588 46294 246612 46350
rect 246668 46294 246736 46350
rect 246792 46294 246860 46350
rect 246916 46294 246984 46350
rect 247040 46294 247064 46350
rect 246588 46226 247064 46294
rect 246588 46170 246612 46226
rect 246668 46170 246736 46226
rect 246792 46170 246860 46226
rect 246916 46170 246984 46226
rect 247040 46170 247064 46226
rect 246588 46102 247064 46170
rect 246588 46046 246612 46102
rect 246668 46046 246736 46102
rect 246792 46046 246860 46102
rect 246916 46046 246984 46102
rect 247040 46046 247064 46102
rect 246588 45978 247064 46046
rect 246588 45922 246612 45978
rect 246668 45922 246736 45978
rect 246792 45922 246860 45978
rect 246916 45922 246984 45978
rect 247040 45922 247064 45978
rect 246588 45888 247064 45922
rect 247772 4676 247828 291452
rect 249228 285684 249284 285694
rect 248768 202350 249088 202384
rect 248768 202294 248838 202350
rect 248894 202294 248962 202350
rect 249018 202294 249088 202350
rect 248768 202226 249088 202294
rect 248768 202170 248838 202226
rect 248894 202170 248962 202226
rect 249018 202170 249088 202226
rect 248768 202102 249088 202170
rect 248768 202046 248838 202102
rect 248894 202046 248962 202102
rect 249018 202046 249088 202102
rect 248768 201978 249088 202046
rect 248768 201922 248838 201978
rect 248894 201922 248962 201978
rect 249018 201922 249088 201978
rect 248768 201888 249088 201922
rect 248768 184350 249088 184384
rect 248768 184294 248838 184350
rect 248894 184294 248962 184350
rect 249018 184294 249088 184350
rect 248768 184226 249088 184294
rect 248768 184170 248838 184226
rect 248894 184170 248962 184226
rect 249018 184170 249088 184226
rect 248768 184102 249088 184170
rect 248768 184046 248838 184102
rect 248894 184046 248962 184102
rect 249018 184046 249088 184102
rect 248768 183978 249088 184046
rect 248768 183922 248838 183978
rect 248894 183922 248962 183978
rect 249018 183922 249088 183978
rect 248768 183888 249088 183922
rect 248768 166350 249088 166384
rect 248768 166294 248838 166350
rect 248894 166294 248962 166350
rect 249018 166294 249088 166350
rect 248768 166226 249088 166294
rect 248768 166170 248838 166226
rect 248894 166170 248962 166226
rect 249018 166170 249088 166226
rect 248768 166102 249088 166170
rect 248768 166046 248838 166102
rect 248894 166046 248962 166102
rect 249018 166046 249088 166102
rect 248768 165978 249088 166046
rect 248768 165922 248838 165978
rect 248894 165922 248962 165978
rect 249018 165922 249088 165978
rect 248768 165888 249088 165922
rect 249228 39508 249284 285628
rect 249228 39442 249284 39452
rect 251178 274350 251798 291922
rect 254898 298350 255518 299890
rect 270508 298788 270564 298798
rect 254898 298294 254994 298350
rect 255050 298294 255118 298350
rect 255174 298294 255242 298350
rect 255298 298294 255366 298350
rect 255422 298294 255518 298350
rect 254898 298226 255518 298294
rect 254898 298170 254994 298226
rect 255050 298170 255118 298226
rect 255174 298170 255242 298226
rect 255298 298170 255366 298226
rect 255422 298170 255518 298226
rect 254898 298102 255518 298170
rect 254898 298046 254994 298102
rect 255050 298046 255118 298102
rect 255174 298046 255242 298102
rect 255298 298046 255366 298102
rect 255422 298046 255518 298102
rect 254898 297978 255518 298046
rect 254898 297922 254994 297978
rect 255050 297922 255118 297978
rect 255174 297922 255242 297978
rect 255298 297922 255366 297978
rect 255422 297922 255518 297978
rect 251178 274294 251274 274350
rect 251330 274294 251398 274350
rect 251454 274294 251522 274350
rect 251578 274294 251646 274350
rect 251702 274294 251798 274350
rect 251178 274226 251798 274294
rect 251178 274170 251274 274226
rect 251330 274170 251398 274226
rect 251454 274170 251522 274226
rect 251578 274170 251646 274226
rect 251702 274170 251798 274226
rect 251178 274102 251798 274170
rect 251178 274046 251274 274102
rect 251330 274046 251398 274102
rect 251454 274046 251522 274102
rect 251578 274046 251646 274102
rect 251702 274046 251798 274102
rect 251178 273978 251798 274046
rect 251178 273922 251274 273978
rect 251330 273922 251398 273978
rect 251454 273922 251522 273978
rect 251578 273922 251646 273978
rect 251702 273922 251798 273978
rect 251178 256350 251798 273922
rect 251178 256294 251274 256350
rect 251330 256294 251398 256350
rect 251454 256294 251522 256350
rect 251578 256294 251646 256350
rect 251702 256294 251798 256350
rect 251178 256226 251798 256294
rect 251178 256170 251274 256226
rect 251330 256170 251398 256226
rect 251454 256170 251522 256226
rect 251578 256170 251646 256226
rect 251702 256170 251798 256226
rect 251178 256102 251798 256170
rect 251178 256046 251274 256102
rect 251330 256046 251398 256102
rect 251454 256046 251522 256102
rect 251578 256046 251646 256102
rect 251702 256046 251798 256102
rect 251178 255978 251798 256046
rect 251178 255922 251274 255978
rect 251330 255922 251398 255978
rect 251454 255922 251522 255978
rect 251578 255922 251646 255978
rect 251702 255922 251798 255978
rect 251178 238350 251798 255922
rect 251178 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 251798 238350
rect 251178 238226 251798 238294
rect 251178 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 251798 238226
rect 251178 238102 251798 238170
rect 251178 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 251798 238102
rect 251178 237978 251798 238046
rect 251178 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 251798 237978
rect 251178 220350 251798 237922
rect 251178 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 251798 220350
rect 251178 220226 251798 220294
rect 251178 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 251798 220226
rect 251178 220102 251798 220170
rect 251178 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 251798 220102
rect 251178 219978 251798 220046
rect 251178 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 251798 219978
rect 251178 202350 251798 219922
rect 251178 202294 251274 202350
rect 251330 202294 251398 202350
rect 251454 202294 251522 202350
rect 251578 202294 251646 202350
rect 251702 202294 251798 202350
rect 251178 202226 251798 202294
rect 251178 202170 251274 202226
rect 251330 202170 251398 202226
rect 251454 202170 251522 202226
rect 251578 202170 251646 202226
rect 251702 202170 251798 202226
rect 251178 202102 251798 202170
rect 251178 202046 251274 202102
rect 251330 202046 251398 202102
rect 251454 202046 251522 202102
rect 251578 202046 251646 202102
rect 251702 202046 251798 202102
rect 251178 201978 251798 202046
rect 251178 201922 251274 201978
rect 251330 201922 251398 201978
rect 251454 201922 251522 201978
rect 251578 201922 251646 201978
rect 251702 201922 251798 201978
rect 251178 184350 251798 201922
rect 251178 184294 251274 184350
rect 251330 184294 251398 184350
rect 251454 184294 251522 184350
rect 251578 184294 251646 184350
rect 251702 184294 251798 184350
rect 251178 184226 251798 184294
rect 251178 184170 251274 184226
rect 251330 184170 251398 184226
rect 251454 184170 251522 184226
rect 251578 184170 251646 184226
rect 251702 184170 251798 184226
rect 251178 184102 251798 184170
rect 251178 184046 251274 184102
rect 251330 184046 251398 184102
rect 251454 184046 251522 184102
rect 251578 184046 251646 184102
rect 251702 184046 251798 184102
rect 251178 183978 251798 184046
rect 251178 183922 251274 183978
rect 251330 183922 251398 183978
rect 251454 183922 251522 183978
rect 251578 183922 251646 183978
rect 251702 183922 251798 183978
rect 251178 166350 251798 183922
rect 251178 166294 251274 166350
rect 251330 166294 251398 166350
rect 251454 166294 251522 166350
rect 251578 166294 251646 166350
rect 251702 166294 251798 166350
rect 251178 166226 251798 166294
rect 251178 166170 251274 166226
rect 251330 166170 251398 166226
rect 251454 166170 251522 166226
rect 251578 166170 251646 166226
rect 251702 166170 251798 166226
rect 251178 166102 251798 166170
rect 251178 166046 251274 166102
rect 251330 166046 251398 166102
rect 251454 166046 251522 166102
rect 251578 166046 251646 166102
rect 251702 166046 251798 166102
rect 251178 165978 251798 166046
rect 251178 165922 251274 165978
rect 251330 165922 251398 165978
rect 251454 165922 251522 165978
rect 251578 165922 251646 165978
rect 251702 165922 251798 165978
rect 251178 148350 251798 165922
rect 251178 148294 251274 148350
rect 251330 148294 251398 148350
rect 251454 148294 251522 148350
rect 251578 148294 251646 148350
rect 251702 148294 251798 148350
rect 251178 148226 251798 148294
rect 251178 148170 251274 148226
rect 251330 148170 251398 148226
rect 251454 148170 251522 148226
rect 251578 148170 251646 148226
rect 251702 148170 251798 148226
rect 251178 148102 251798 148170
rect 251178 148046 251274 148102
rect 251330 148046 251398 148102
rect 251454 148046 251522 148102
rect 251578 148046 251646 148102
rect 251702 148046 251798 148102
rect 251178 147978 251798 148046
rect 251178 147922 251274 147978
rect 251330 147922 251398 147978
rect 251454 147922 251522 147978
rect 251578 147922 251646 147978
rect 251702 147922 251798 147978
rect 251178 130350 251798 147922
rect 251178 130294 251274 130350
rect 251330 130294 251398 130350
rect 251454 130294 251522 130350
rect 251578 130294 251646 130350
rect 251702 130294 251798 130350
rect 251178 130226 251798 130294
rect 251178 130170 251274 130226
rect 251330 130170 251398 130226
rect 251454 130170 251522 130226
rect 251578 130170 251646 130226
rect 251702 130170 251798 130226
rect 251178 130102 251798 130170
rect 251178 130046 251274 130102
rect 251330 130046 251398 130102
rect 251454 130046 251522 130102
rect 251578 130046 251646 130102
rect 251702 130046 251798 130102
rect 251178 129978 251798 130046
rect 251178 129922 251274 129978
rect 251330 129922 251398 129978
rect 251454 129922 251522 129978
rect 251578 129922 251646 129978
rect 251702 129922 251798 129978
rect 251178 112350 251798 129922
rect 251178 112294 251274 112350
rect 251330 112294 251398 112350
rect 251454 112294 251522 112350
rect 251578 112294 251646 112350
rect 251702 112294 251798 112350
rect 251178 112226 251798 112294
rect 251178 112170 251274 112226
rect 251330 112170 251398 112226
rect 251454 112170 251522 112226
rect 251578 112170 251646 112226
rect 251702 112170 251798 112226
rect 251178 112102 251798 112170
rect 251178 112046 251274 112102
rect 251330 112046 251398 112102
rect 251454 112046 251522 112102
rect 251578 112046 251646 112102
rect 251702 112046 251798 112102
rect 251178 111978 251798 112046
rect 251178 111922 251274 111978
rect 251330 111922 251398 111978
rect 251454 111922 251522 111978
rect 251578 111922 251646 111978
rect 251702 111922 251798 111978
rect 251178 94350 251798 111922
rect 251178 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 251798 94350
rect 251178 94226 251798 94294
rect 251178 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 251798 94226
rect 251178 94102 251798 94170
rect 251178 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 251798 94102
rect 251178 93978 251798 94046
rect 251178 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 251798 93978
rect 251178 76350 251798 93922
rect 251178 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 251798 76350
rect 251178 76226 251798 76294
rect 251178 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 251798 76226
rect 251178 76102 251798 76170
rect 251178 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 251798 76102
rect 251178 75978 251798 76046
rect 251178 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 251798 75978
rect 251178 58350 251798 75922
rect 251178 58294 251274 58350
rect 251330 58294 251398 58350
rect 251454 58294 251522 58350
rect 251578 58294 251646 58350
rect 251702 58294 251798 58350
rect 251178 58226 251798 58294
rect 251178 58170 251274 58226
rect 251330 58170 251398 58226
rect 251454 58170 251522 58226
rect 251578 58170 251646 58226
rect 251702 58170 251798 58226
rect 251178 58102 251798 58170
rect 251178 58046 251274 58102
rect 251330 58046 251398 58102
rect 251454 58046 251522 58102
rect 251578 58046 251646 58102
rect 251702 58046 251798 58102
rect 251178 57978 251798 58046
rect 251178 57922 251274 57978
rect 251330 57922 251398 57978
rect 251454 57922 251522 57978
rect 251578 57922 251646 57978
rect 251702 57922 251798 57978
rect 251178 40350 251798 57922
rect 251178 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 251798 40350
rect 251178 40226 251798 40294
rect 251178 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 251798 40226
rect 251178 40102 251798 40170
rect 251178 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 251798 40102
rect 251178 39978 251798 40046
rect 251178 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 251798 39978
rect 247772 4610 247828 4620
rect 251178 22350 251798 39922
rect 251178 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 251798 22350
rect 251178 22226 251798 22294
rect 251178 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 251798 22226
rect 251178 22102 251798 22170
rect 251178 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 251798 22102
rect 251178 21978 251798 22046
rect 251178 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 251798 21978
rect 245196 4162 245252 4172
rect 251178 4350 251798 21922
rect 252028 285796 252084 285806
rect 252028 7588 252084 285740
rect 252140 285684 252196 285694
rect 252140 37940 252196 285628
rect 252140 37874 252196 37884
rect 254898 280350 255518 297922
rect 264128 298350 264448 298384
rect 264128 298294 264198 298350
rect 264254 298294 264322 298350
rect 264378 298294 264448 298350
rect 264128 298226 264448 298294
rect 264128 298170 264198 298226
rect 264254 298170 264322 298226
rect 264378 298170 264448 298226
rect 264128 298102 264448 298170
rect 264128 298046 264198 298102
rect 264254 298046 264322 298102
rect 264378 298046 264448 298102
rect 264128 297978 264448 298046
rect 264128 297922 264198 297978
rect 264254 297922 264322 297978
rect 264378 297922 264448 297978
rect 264128 297888 264448 297922
rect 269388 297444 269444 297454
rect 258748 286468 258804 286478
rect 255724 286356 255780 286366
rect 254898 280294 254994 280350
rect 255050 280294 255118 280350
rect 255174 280294 255242 280350
rect 255298 280294 255366 280350
rect 255422 280294 255518 280350
rect 254898 280226 255518 280294
rect 254898 280170 254994 280226
rect 255050 280170 255118 280226
rect 255174 280170 255242 280226
rect 255298 280170 255366 280226
rect 255422 280170 255518 280226
rect 254898 280102 255518 280170
rect 254898 280046 254994 280102
rect 255050 280046 255118 280102
rect 255174 280046 255242 280102
rect 255298 280046 255366 280102
rect 255422 280046 255518 280102
rect 254898 279978 255518 280046
rect 254898 279922 254994 279978
rect 255050 279922 255118 279978
rect 255174 279922 255242 279978
rect 255298 279922 255366 279978
rect 255422 279922 255518 279978
rect 254898 262350 255518 279922
rect 254898 262294 254994 262350
rect 255050 262294 255118 262350
rect 255174 262294 255242 262350
rect 255298 262294 255366 262350
rect 255422 262294 255518 262350
rect 254898 262226 255518 262294
rect 254898 262170 254994 262226
rect 255050 262170 255118 262226
rect 255174 262170 255242 262226
rect 255298 262170 255366 262226
rect 255422 262170 255518 262226
rect 254898 262102 255518 262170
rect 254898 262046 254994 262102
rect 255050 262046 255118 262102
rect 255174 262046 255242 262102
rect 255298 262046 255366 262102
rect 255422 262046 255518 262102
rect 254898 261978 255518 262046
rect 254898 261922 254994 261978
rect 255050 261922 255118 261978
rect 255174 261922 255242 261978
rect 255298 261922 255366 261978
rect 255422 261922 255518 261978
rect 254898 244350 255518 261922
rect 254898 244294 254994 244350
rect 255050 244294 255118 244350
rect 255174 244294 255242 244350
rect 255298 244294 255366 244350
rect 255422 244294 255518 244350
rect 254898 244226 255518 244294
rect 254898 244170 254994 244226
rect 255050 244170 255118 244226
rect 255174 244170 255242 244226
rect 255298 244170 255366 244226
rect 255422 244170 255518 244226
rect 254898 244102 255518 244170
rect 254898 244046 254994 244102
rect 255050 244046 255118 244102
rect 255174 244046 255242 244102
rect 255298 244046 255366 244102
rect 255422 244046 255518 244102
rect 254898 243978 255518 244046
rect 254898 243922 254994 243978
rect 255050 243922 255118 243978
rect 255174 243922 255242 243978
rect 255298 243922 255366 243978
rect 255422 243922 255518 243978
rect 254898 226350 255518 243922
rect 254898 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 255518 226350
rect 254898 226226 255518 226294
rect 254898 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 255518 226226
rect 254898 226102 255518 226170
rect 254898 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 255518 226102
rect 254898 225978 255518 226046
rect 254898 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 255518 225978
rect 254898 208350 255518 225922
rect 254898 208294 254994 208350
rect 255050 208294 255118 208350
rect 255174 208294 255242 208350
rect 255298 208294 255366 208350
rect 255422 208294 255518 208350
rect 254898 208226 255518 208294
rect 254898 208170 254994 208226
rect 255050 208170 255118 208226
rect 255174 208170 255242 208226
rect 255298 208170 255366 208226
rect 255422 208170 255518 208226
rect 254898 208102 255518 208170
rect 254898 208046 254994 208102
rect 255050 208046 255118 208102
rect 255174 208046 255242 208102
rect 255298 208046 255366 208102
rect 255422 208046 255518 208102
rect 254898 207978 255518 208046
rect 254898 207922 254994 207978
rect 255050 207922 255118 207978
rect 255174 207922 255242 207978
rect 255298 207922 255366 207978
rect 255422 207922 255518 207978
rect 254898 190350 255518 207922
rect 254898 190294 254994 190350
rect 255050 190294 255118 190350
rect 255174 190294 255242 190350
rect 255298 190294 255366 190350
rect 255422 190294 255518 190350
rect 254898 190226 255518 190294
rect 254898 190170 254994 190226
rect 255050 190170 255118 190226
rect 255174 190170 255242 190226
rect 255298 190170 255366 190226
rect 255422 190170 255518 190226
rect 254898 190102 255518 190170
rect 254898 190046 254994 190102
rect 255050 190046 255118 190102
rect 255174 190046 255242 190102
rect 255298 190046 255366 190102
rect 255422 190046 255518 190102
rect 254898 189978 255518 190046
rect 254898 189922 254994 189978
rect 255050 189922 255118 189978
rect 255174 189922 255242 189978
rect 255298 189922 255366 189978
rect 255422 189922 255518 189978
rect 254898 172350 255518 189922
rect 254898 172294 254994 172350
rect 255050 172294 255118 172350
rect 255174 172294 255242 172350
rect 255298 172294 255366 172350
rect 255422 172294 255518 172350
rect 254898 172226 255518 172294
rect 254898 172170 254994 172226
rect 255050 172170 255118 172226
rect 255174 172170 255242 172226
rect 255298 172170 255366 172226
rect 255422 172170 255518 172226
rect 254898 172102 255518 172170
rect 254898 172046 254994 172102
rect 255050 172046 255118 172102
rect 255174 172046 255242 172102
rect 255298 172046 255366 172102
rect 255422 172046 255518 172102
rect 254898 171978 255518 172046
rect 254898 171922 254994 171978
rect 255050 171922 255118 171978
rect 255174 171922 255242 171978
rect 255298 171922 255366 171978
rect 255422 171922 255518 171978
rect 254898 154350 255518 171922
rect 254898 154294 254994 154350
rect 255050 154294 255118 154350
rect 255174 154294 255242 154350
rect 255298 154294 255366 154350
rect 255422 154294 255518 154350
rect 254898 154226 255518 154294
rect 254898 154170 254994 154226
rect 255050 154170 255118 154226
rect 255174 154170 255242 154226
rect 255298 154170 255366 154226
rect 255422 154170 255518 154226
rect 254898 154102 255518 154170
rect 254898 154046 254994 154102
rect 255050 154046 255118 154102
rect 255174 154046 255242 154102
rect 255298 154046 255366 154102
rect 255422 154046 255518 154102
rect 254898 153978 255518 154046
rect 254898 153922 254994 153978
rect 255050 153922 255118 153978
rect 255174 153922 255242 153978
rect 255298 153922 255366 153978
rect 255422 153922 255518 153978
rect 254898 136350 255518 153922
rect 254898 136294 254994 136350
rect 255050 136294 255118 136350
rect 255174 136294 255242 136350
rect 255298 136294 255366 136350
rect 255422 136294 255518 136350
rect 254898 136226 255518 136294
rect 254898 136170 254994 136226
rect 255050 136170 255118 136226
rect 255174 136170 255242 136226
rect 255298 136170 255366 136226
rect 255422 136170 255518 136226
rect 254898 136102 255518 136170
rect 254898 136046 254994 136102
rect 255050 136046 255118 136102
rect 255174 136046 255242 136102
rect 255298 136046 255366 136102
rect 255422 136046 255518 136102
rect 254898 135978 255518 136046
rect 254898 135922 254994 135978
rect 255050 135922 255118 135978
rect 255174 135922 255242 135978
rect 255298 135922 255366 135978
rect 255422 135922 255518 135978
rect 254898 118350 255518 135922
rect 254898 118294 254994 118350
rect 255050 118294 255118 118350
rect 255174 118294 255242 118350
rect 255298 118294 255366 118350
rect 255422 118294 255518 118350
rect 254898 118226 255518 118294
rect 254898 118170 254994 118226
rect 255050 118170 255118 118226
rect 255174 118170 255242 118226
rect 255298 118170 255366 118226
rect 255422 118170 255518 118226
rect 254898 118102 255518 118170
rect 254898 118046 254994 118102
rect 255050 118046 255118 118102
rect 255174 118046 255242 118102
rect 255298 118046 255366 118102
rect 255422 118046 255518 118102
rect 254898 117978 255518 118046
rect 254898 117922 254994 117978
rect 255050 117922 255118 117978
rect 255174 117922 255242 117978
rect 255298 117922 255366 117978
rect 255422 117922 255518 117978
rect 254898 100350 255518 117922
rect 254898 100294 254994 100350
rect 255050 100294 255118 100350
rect 255174 100294 255242 100350
rect 255298 100294 255366 100350
rect 255422 100294 255518 100350
rect 254898 100226 255518 100294
rect 254898 100170 254994 100226
rect 255050 100170 255118 100226
rect 255174 100170 255242 100226
rect 255298 100170 255366 100226
rect 255422 100170 255518 100226
rect 254898 100102 255518 100170
rect 254898 100046 254994 100102
rect 255050 100046 255118 100102
rect 255174 100046 255242 100102
rect 255298 100046 255366 100102
rect 255422 100046 255518 100102
rect 254898 99978 255518 100046
rect 254898 99922 254994 99978
rect 255050 99922 255118 99978
rect 255174 99922 255242 99978
rect 255298 99922 255366 99978
rect 255422 99922 255518 99978
rect 254898 82350 255518 99922
rect 254898 82294 254994 82350
rect 255050 82294 255118 82350
rect 255174 82294 255242 82350
rect 255298 82294 255366 82350
rect 255422 82294 255518 82350
rect 254898 82226 255518 82294
rect 254898 82170 254994 82226
rect 255050 82170 255118 82226
rect 255174 82170 255242 82226
rect 255298 82170 255366 82226
rect 255422 82170 255518 82226
rect 254898 82102 255518 82170
rect 254898 82046 254994 82102
rect 255050 82046 255118 82102
rect 255174 82046 255242 82102
rect 255298 82046 255366 82102
rect 255422 82046 255518 82102
rect 254898 81978 255518 82046
rect 254898 81922 254994 81978
rect 255050 81922 255118 81978
rect 255174 81922 255242 81978
rect 255298 81922 255366 81978
rect 255422 81922 255518 81978
rect 254898 64350 255518 81922
rect 254898 64294 254994 64350
rect 255050 64294 255118 64350
rect 255174 64294 255242 64350
rect 255298 64294 255366 64350
rect 255422 64294 255518 64350
rect 254898 64226 255518 64294
rect 254898 64170 254994 64226
rect 255050 64170 255118 64226
rect 255174 64170 255242 64226
rect 255298 64170 255366 64226
rect 255422 64170 255518 64226
rect 254898 64102 255518 64170
rect 254898 64046 254994 64102
rect 255050 64046 255118 64102
rect 255174 64046 255242 64102
rect 255298 64046 255366 64102
rect 255422 64046 255518 64102
rect 254898 63978 255518 64046
rect 254898 63922 254994 63978
rect 255050 63922 255118 63978
rect 255174 63922 255242 63978
rect 255298 63922 255366 63978
rect 255422 63922 255518 63978
rect 254898 46350 255518 63922
rect 254898 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 255518 46350
rect 254898 46226 255518 46294
rect 254898 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 255518 46226
rect 254898 46102 255518 46170
rect 254898 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 255518 46102
rect 254898 45978 255518 46046
rect 254898 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 255518 45978
rect 252028 7522 252084 7532
rect 254898 28350 255518 45922
rect 255612 285684 255668 285694
rect 255612 36148 255668 285628
rect 255724 37828 255780 286300
rect 257964 285908 258020 285918
rect 255724 37762 255780 37772
rect 257852 285684 257908 285694
rect 255612 36082 255668 36092
rect 257852 31108 257908 285628
rect 257964 32788 258020 285852
rect 257964 32722 258020 32732
rect 257852 31042 257908 31052
rect 258748 29428 258804 286412
rect 259532 285796 259588 285806
rect 259532 36260 259588 285740
rect 260428 285684 260484 285694
rect 260428 138964 260484 285628
rect 265468 285684 265524 285694
rect 264128 190350 264448 190384
rect 264128 190294 264198 190350
rect 264254 190294 264322 190350
rect 264378 190294 264448 190350
rect 264128 190226 264448 190294
rect 264128 190170 264198 190226
rect 264254 190170 264322 190226
rect 264378 190170 264448 190226
rect 264128 190102 264448 190170
rect 264128 190046 264198 190102
rect 264254 190046 264322 190102
rect 264378 190046 264448 190102
rect 264128 189978 264448 190046
rect 264128 189922 264198 189978
rect 264254 189922 264322 189978
rect 264378 189922 264448 189978
rect 264128 189888 264448 189922
rect 264128 172350 264448 172384
rect 264128 172294 264198 172350
rect 264254 172294 264322 172350
rect 264378 172294 264448 172350
rect 264128 172226 264448 172294
rect 264128 172170 264198 172226
rect 264254 172170 264322 172226
rect 264378 172170 264448 172226
rect 264128 172102 264448 172170
rect 264128 172046 264198 172102
rect 264254 172046 264322 172102
rect 264378 172046 264448 172102
rect 264128 171978 264448 172046
rect 264128 171922 264198 171978
rect 264254 171922 264322 171978
rect 264378 171922 264448 171978
rect 264128 171888 264448 171922
rect 265468 151172 265524 285628
rect 265468 151106 265524 151116
rect 267036 160244 267092 160254
rect 260428 138898 260484 138908
rect 261106 130350 261582 130384
rect 261106 130294 261130 130350
rect 261186 130294 261254 130350
rect 261310 130294 261378 130350
rect 261434 130294 261502 130350
rect 261558 130294 261582 130350
rect 261106 130226 261582 130294
rect 261106 130170 261130 130226
rect 261186 130170 261254 130226
rect 261310 130170 261378 130226
rect 261434 130170 261502 130226
rect 261558 130170 261582 130226
rect 261106 130102 261582 130170
rect 261106 130046 261130 130102
rect 261186 130046 261254 130102
rect 261310 130046 261378 130102
rect 261434 130046 261502 130102
rect 261558 130046 261582 130102
rect 261106 129978 261582 130046
rect 261106 129922 261130 129978
rect 261186 129922 261254 129978
rect 261310 129922 261378 129978
rect 261434 129922 261502 129978
rect 261558 129922 261582 129978
rect 261106 129888 261582 129922
rect 261906 118350 262382 118384
rect 261906 118294 261930 118350
rect 261986 118294 262054 118350
rect 262110 118294 262178 118350
rect 262234 118294 262302 118350
rect 262358 118294 262382 118350
rect 261906 118226 262382 118294
rect 261906 118170 261930 118226
rect 261986 118170 262054 118226
rect 262110 118170 262178 118226
rect 262234 118170 262302 118226
rect 262358 118170 262382 118226
rect 261906 118102 262382 118170
rect 261906 118046 261930 118102
rect 261986 118046 262054 118102
rect 262110 118046 262178 118102
rect 262234 118046 262302 118102
rect 262358 118046 262382 118102
rect 261906 117978 262382 118046
rect 261906 117922 261930 117978
rect 261986 117922 262054 117978
rect 262110 117922 262178 117978
rect 262234 117922 262302 117978
rect 262358 117922 262382 117978
rect 261906 117888 262382 117922
rect 261106 112350 261582 112384
rect 261106 112294 261130 112350
rect 261186 112294 261254 112350
rect 261310 112294 261378 112350
rect 261434 112294 261502 112350
rect 261558 112294 261582 112350
rect 261106 112226 261582 112294
rect 261106 112170 261130 112226
rect 261186 112170 261254 112226
rect 261310 112170 261378 112226
rect 261434 112170 261502 112226
rect 261558 112170 261582 112226
rect 261106 112102 261582 112170
rect 261106 112046 261130 112102
rect 261186 112046 261254 112102
rect 261310 112046 261378 112102
rect 261434 112046 261502 112102
rect 261558 112046 261582 112102
rect 261106 111978 261582 112046
rect 261106 111922 261130 111978
rect 261186 111922 261254 111978
rect 261310 111922 261378 111978
rect 261434 111922 261502 111978
rect 261558 111922 261582 111978
rect 261106 111888 261582 111922
rect 261906 100350 262382 100384
rect 261906 100294 261930 100350
rect 261986 100294 262054 100350
rect 262110 100294 262178 100350
rect 262234 100294 262302 100350
rect 262358 100294 262382 100350
rect 261906 100226 262382 100294
rect 261906 100170 261930 100226
rect 261986 100170 262054 100226
rect 262110 100170 262178 100226
rect 262234 100170 262302 100226
rect 262358 100170 262382 100226
rect 261906 100102 262382 100170
rect 261906 100046 261930 100102
rect 261986 100046 262054 100102
rect 262110 100046 262178 100102
rect 262234 100046 262302 100102
rect 262358 100046 262382 100102
rect 261906 99978 262382 100046
rect 261906 99922 261930 99978
rect 261986 99922 262054 99978
rect 262110 99922 262178 99978
rect 262234 99922 262302 99978
rect 262358 99922 262382 99978
rect 261906 99888 262382 99922
rect 261106 94350 261582 94384
rect 261106 94294 261130 94350
rect 261186 94294 261254 94350
rect 261310 94294 261378 94350
rect 261434 94294 261502 94350
rect 261558 94294 261582 94350
rect 261106 94226 261582 94294
rect 261106 94170 261130 94226
rect 261186 94170 261254 94226
rect 261310 94170 261378 94226
rect 261434 94170 261502 94226
rect 261558 94170 261582 94226
rect 261106 94102 261582 94170
rect 261106 94046 261130 94102
rect 261186 94046 261254 94102
rect 261310 94046 261378 94102
rect 261434 94046 261502 94102
rect 261558 94046 261582 94102
rect 261106 93978 261582 94046
rect 261106 93922 261130 93978
rect 261186 93922 261254 93978
rect 261310 93922 261378 93978
rect 261434 93922 261502 93978
rect 261558 93922 261582 93978
rect 261106 93888 261582 93922
rect 261906 82350 262382 82384
rect 261906 82294 261930 82350
rect 261986 82294 262054 82350
rect 262110 82294 262178 82350
rect 262234 82294 262302 82350
rect 262358 82294 262382 82350
rect 261906 82226 262382 82294
rect 261906 82170 261930 82226
rect 261986 82170 262054 82226
rect 262110 82170 262178 82226
rect 262234 82170 262302 82226
rect 262358 82170 262382 82226
rect 261906 82102 262382 82170
rect 261906 82046 261930 82102
rect 261986 82046 262054 82102
rect 262110 82046 262178 82102
rect 262234 82046 262302 82102
rect 262358 82046 262382 82102
rect 261906 81978 262382 82046
rect 261906 81922 261930 81978
rect 261986 81922 262054 81978
rect 262110 81922 262178 81978
rect 262234 81922 262302 81978
rect 262358 81922 262382 81978
rect 261906 81888 262382 81922
rect 261106 76350 261582 76384
rect 261106 76294 261130 76350
rect 261186 76294 261254 76350
rect 261310 76294 261378 76350
rect 261434 76294 261502 76350
rect 261558 76294 261582 76350
rect 261106 76226 261582 76294
rect 261106 76170 261130 76226
rect 261186 76170 261254 76226
rect 261310 76170 261378 76226
rect 261434 76170 261502 76226
rect 261558 76170 261582 76226
rect 261106 76102 261582 76170
rect 261106 76046 261130 76102
rect 261186 76046 261254 76102
rect 261310 76046 261378 76102
rect 261434 76046 261502 76102
rect 261558 76046 261582 76102
rect 261106 75978 261582 76046
rect 261106 75922 261130 75978
rect 261186 75922 261254 75978
rect 261310 75922 261378 75978
rect 261434 75922 261502 75978
rect 261558 75922 261582 75978
rect 261106 75888 261582 75922
rect 261906 64350 262382 64384
rect 261906 64294 261930 64350
rect 261986 64294 262054 64350
rect 262110 64294 262178 64350
rect 262234 64294 262302 64350
rect 262358 64294 262382 64350
rect 261906 64226 262382 64294
rect 261906 64170 261930 64226
rect 261986 64170 262054 64226
rect 262110 64170 262178 64226
rect 262234 64170 262302 64226
rect 262358 64170 262382 64226
rect 261906 64102 262382 64170
rect 261906 64046 261930 64102
rect 261986 64046 262054 64102
rect 262110 64046 262178 64102
rect 262234 64046 262302 64102
rect 262358 64046 262382 64102
rect 261906 63978 262382 64046
rect 261906 63922 261930 63978
rect 261986 63922 262054 63978
rect 262110 63922 262178 63978
rect 262234 63922 262302 63978
rect 262358 63922 262382 63978
rect 261906 63888 262382 63922
rect 261106 58350 261582 58384
rect 261106 58294 261130 58350
rect 261186 58294 261254 58350
rect 261310 58294 261378 58350
rect 261434 58294 261502 58350
rect 261558 58294 261582 58350
rect 261106 58226 261582 58294
rect 261106 58170 261130 58226
rect 261186 58170 261254 58226
rect 261310 58170 261378 58226
rect 261434 58170 261502 58226
rect 261558 58170 261582 58226
rect 261106 58102 261582 58170
rect 261106 58046 261130 58102
rect 261186 58046 261254 58102
rect 261310 58046 261378 58102
rect 261434 58046 261502 58102
rect 261558 58046 261582 58102
rect 261106 57978 261582 58046
rect 261106 57922 261130 57978
rect 261186 57922 261254 57978
rect 261310 57922 261378 57978
rect 261434 57922 261502 57978
rect 261558 57922 261582 57978
rect 261106 57888 261582 57922
rect 261906 46350 262382 46384
rect 261906 46294 261930 46350
rect 261986 46294 262054 46350
rect 262110 46294 262178 46350
rect 262234 46294 262302 46350
rect 262358 46294 262382 46350
rect 261906 46226 262382 46294
rect 261906 46170 261930 46226
rect 261986 46170 262054 46226
rect 262110 46170 262178 46226
rect 262234 46170 262302 46226
rect 262358 46170 262382 46226
rect 261906 46102 262382 46170
rect 261906 46046 261930 46102
rect 261986 46046 262054 46102
rect 262110 46046 262178 46102
rect 262234 46046 262302 46102
rect 262358 46046 262382 46102
rect 261906 45978 262382 46046
rect 261906 45922 261930 45978
rect 261986 45922 262054 45978
rect 262110 45922 262178 45978
rect 262234 45922 262302 45978
rect 262358 45922 262382 45978
rect 261906 45888 262382 45922
rect 259532 36194 259588 36204
rect 258748 29362 258804 29372
rect 254898 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 255518 28350
rect 254898 28226 255518 28294
rect 254898 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 255518 28226
rect 254898 28102 255518 28170
rect 254898 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 255518 28102
rect 254898 27978 255518 28046
rect 254898 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 255518 27978
rect 254898 10350 255518 27922
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 233436 4050 233492 4060
rect 251178 4102 251798 4170
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 251178 -160 251798 3922
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 -1120 255518 9922
rect 267036 4340 267092 160188
rect 269388 5908 269444 297388
rect 270508 6020 270564 298732
rect 272188 148820 272244 310828
rect 272188 148754 272244 148764
rect 273868 308196 273924 308206
rect 273868 14308 273924 308140
rect 274652 291620 274708 317582
rect 277676 312228 277732 312238
rect 276332 307558 276388 307568
rect 276332 291732 276388 307502
rect 276332 291666 276388 291676
rect 274652 291554 274708 291564
rect 277676 20188 277732 312172
rect 278236 291844 278292 376442
rect 279692 337618 279748 429100
rect 281372 427258 281428 427268
rect 281372 345718 281428 427202
rect 281372 345652 281428 345662
rect 281898 418350 282518 435922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 568350 286238 585922
rect 285618 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 286238 568350
rect 285618 568226 286238 568294
rect 285618 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 286238 568226
rect 285618 568102 286238 568170
rect 285618 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 286238 568102
rect 285618 567978 286238 568046
rect 285618 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 286238 567978
rect 285618 550350 286238 567922
rect 285618 550294 285714 550350
rect 285770 550294 285838 550350
rect 285894 550294 285962 550350
rect 286018 550294 286086 550350
rect 286142 550294 286238 550350
rect 285618 550226 286238 550294
rect 285618 550170 285714 550226
rect 285770 550170 285838 550226
rect 285894 550170 285962 550226
rect 286018 550170 286086 550226
rect 286142 550170 286238 550226
rect 285618 550102 286238 550170
rect 285618 550046 285714 550102
rect 285770 550046 285838 550102
rect 285894 550046 285962 550102
rect 286018 550046 286086 550102
rect 286142 550046 286238 550102
rect 285618 549978 286238 550046
rect 285618 549922 285714 549978
rect 285770 549922 285838 549978
rect 285894 549922 285962 549978
rect 286018 549922 286086 549978
rect 286142 549922 286238 549978
rect 285618 532350 286238 549922
rect 285618 532294 285714 532350
rect 285770 532294 285838 532350
rect 285894 532294 285962 532350
rect 286018 532294 286086 532350
rect 286142 532294 286238 532350
rect 285618 532226 286238 532294
rect 285618 532170 285714 532226
rect 285770 532170 285838 532226
rect 285894 532170 285962 532226
rect 286018 532170 286086 532226
rect 286142 532170 286238 532226
rect 285618 532102 286238 532170
rect 285618 532046 285714 532102
rect 285770 532046 285838 532102
rect 285894 532046 285962 532102
rect 286018 532046 286086 532102
rect 286142 532046 286238 532102
rect 285618 531978 286238 532046
rect 285618 531922 285714 531978
rect 285770 531922 285838 531978
rect 285894 531922 285962 531978
rect 286018 531922 286086 531978
rect 286142 531922 286238 531978
rect 285618 514350 286238 531922
rect 285618 514294 285714 514350
rect 285770 514294 285838 514350
rect 285894 514294 285962 514350
rect 286018 514294 286086 514350
rect 286142 514294 286238 514350
rect 285618 514226 286238 514294
rect 285618 514170 285714 514226
rect 285770 514170 285838 514226
rect 285894 514170 285962 514226
rect 286018 514170 286086 514226
rect 286142 514170 286238 514226
rect 285618 514102 286238 514170
rect 285618 514046 285714 514102
rect 285770 514046 285838 514102
rect 285894 514046 285962 514102
rect 286018 514046 286086 514102
rect 286142 514046 286238 514102
rect 285618 513978 286238 514046
rect 285618 513922 285714 513978
rect 285770 513922 285838 513978
rect 285894 513922 285962 513978
rect 286018 513922 286086 513978
rect 286142 513922 286238 513978
rect 285618 496350 286238 513922
rect 285618 496294 285714 496350
rect 285770 496294 285838 496350
rect 285894 496294 285962 496350
rect 286018 496294 286086 496350
rect 286142 496294 286238 496350
rect 285618 496226 286238 496294
rect 285618 496170 285714 496226
rect 285770 496170 285838 496226
rect 285894 496170 285962 496226
rect 286018 496170 286086 496226
rect 286142 496170 286238 496226
rect 285618 496102 286238 496170
rect 285618 496046 285714 496102
rect 285770 496046 285838 496102
rect 285894 496046 285962 496102
rect 286018 496046 286086 496102
rect 286142 496046 286238 496102
rect 285618 495978 286238 496046
rect 285618 495922 285714 495978
rect 285770 495922 285838 495978
rect 285894 495922 285962 495978
rect 286018 495922 286086 495978
rect 286142 495922 286238 495978
rect 285618 478350 286238 495922
rect 285618 478294 285714 478350
rect 285770 478294 285838 478350
rect 285894 478294 285962 478350
rect 286018 478294 286086 478350
rect 286142 478294 286238 478350
rect 285618 478226 286238 478294
rect 285618 478170 285714 478226
rect 285770 478170 285838 478226
rect 285894 478170 285962 478226
rect 286018 478170 286086 478226
rect 286142 478170 286238 478226
rect 285618 478102 286238 478170
rect 285618 478046 285714 478102
rect 285770 478046 285838 478102
rect 285894 478046 285962 478102
rect 286018 478046 286086 478102
rect 286142 478046 286238 478102
rect 285618 477978 286238 478046
rect 285618 477922 285714 477978
rect 285770 477922 285838 477978
rect 285894 477922 285962 477978
rect 286018 477922 286086 477978
rect 286142 477922 286238 477978
rect 285618 460350 286238 477922
rect 285618 460294 285714 460350
rect 285770 460294 285838 460350
rect 285894 460294 285962 460350
rect 286018 460294 286086 460350
rect 286142 460294 286238 460350
rect 285618 460226 286238 460294
rect 285618 460170 285714 460226
rect 285770 460170 285838 460226
rect 285894 460170 285962 460226
rect 286018 460170 286086 460226
rect 286142 460170 286238 460226
rect 285618 460102 286238 460170
rect 285618 460046 285714 460102
rect 285770 460046 285838 460102
rect 285894 460046 285962 460102
rect 286018 460046 286086 460102
rect 286142 460046 286238 460102
rect 285618 459978 286238 460046
rect 285618 459922 285714 459978
rect 285770 459922 285838 459978
rect 285894 459922 285962 459978
rect 286018 459922 286086 459978
rect 286142 459922 286238 459978
rect 285618 442350 286238 459922
rect 285618 442294 285714 442350
rect 285770 442294 285838 442350
rect 285894 442294 285962 442350
rect 286018 442294 286086 442350
rect 286142 442294 286238 442350
rect 285618 442226 286238 442294
rect 285618 442170 285714 442226
rect 285770 442170 285838 442226
rect 285894 442170 285962 442226
rect 286018 442170 286086 442226
rect 286142 442170 286238 442226
rect 285618 442102 286238 442170
rect 285618 442046 285714 442102
rect 285770 442046 285838 442102
rect 285894 442046 285962 442102
rect 286018 442046 286086 442102
rect 286142 442046 286238 442102
rect 285618 441978 286238 442046
rect 285618 441922 285714 441978
rect 285770 441922 285838 441978
rect 285894 441922 285962 441978
rect 286018 441922 286086 441978
rect 286142 441922 286238 441978
rect 284844 429418 284900 429428
rect 281898 418294 281994 418350
rect 282050 418294 282118 418350
rect 282174 418294 282242 418350
rect 282298 418294 282366 418350
rect 282422 418294 282518 418350
rect 281898 418226 282518 418294
rect 281898 418170 281994 418226
rect 282050 418170 282118 418226
rect 282174 418170 282242 418226
rect 282298 418170 282366 418226
rect 282422 418170 282518 418226
rect 281898 418102 282518 418170
rect 281898 418046 281994 418102
rect 282050 418046 282118 418102
rect 282174 418046 282242 418102
rect 282298 418046 282366 418102
rect 282422 418046 282518 418102
rect 281898 417978 282518 418046
rect 281898 417922 281994 417978
rect 282050 417922 282118 417978
rect 282174 417922 282242 417978
rect 282298 417922 282366 417978
rect 282422 417922 282518 417978
rect 281898 400350 282518 417922
rect 281898 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 282518 400350
rect 281898 400226 282518 400294
rect 281898 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 282518 400226
rect 281898 400102 282518 400170
rect 281898 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 282518 400102
rect 281898 399978 282518 400046
rect 281898 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 282518 399978
rect 281898 382350 282518 399922
rect 281898 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 282518 382350
rect 281898 382226 282518 382294
rect 281898 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 282518 382226
rect 281898 382102 282518 382170
rect 281898 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 282518 382102
rect 281898 381978 282518 382046
rect 281898 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 282518 381978
rect 281898 364350 282518 381922
rect 281898 364294 281994 364350
rect 282050 364294 282118 364350
rect 282174 364294 282242 364350
rect 282298 364294 282366 364350
rect 282422 364294 282518 364350
rect 281898 364226 282518 364294
rect 281898 364170 281994 364226
rect 282050 364170 282118 364226
rect 282174 364170 282242 364226
rect 282298 364170 282366 364226
rect 282422 364170 282518 364226
rect 281898 364102 282518 364170
rect 281898 364046 281994 364102
rect 282050 364046 282118 364102
rect 282174 364046 282242 364102
rect 282298 364046 282366 364102
rect 282422 364046 282518 364102
rect 281898 363978 282518 364046
rect 281898 363922 281994 363978
rect 282050 363922 282118 363978
rect 282174 363922 282242 363978
rect 282298 363922 282366 363978
rect 282422 363922 282518 363978
rect 281898 346350 282518 363922
rect 281898 346294 281994 346350
rect 282050 346294 282118 346350
rect 282174 346294 282242 346350
rect 282298 346294 282366 346350
rect 282422 346294 282518 346350
rect 281898 346226 282518 346294
rect 281898 346170 281994 346226
rect 282050 346170 282118 346226
rect 282174 346170 282242 346226
rect 282298 346170 282366 346226
rect 282422 346170 282518 346226
rect 281898 346102 282518 346170
rect 281898 346046 281994 346102
rect 282050 346046 282118 346102
rect 282174 346046 282242 346102
rect 282298 346046 282366 346102
rect 282422 346046 282518 346102
rect 281898 345978 282518 346046
rect 281898 345922 281994 345978
rect 282050 345922 282118 345978
rect 282174 345922 282242 345978
rect 282298 345922 282366 345978
rect 282422 345922 282518 345978
rect 279692 337552 279748 337562
rect 281898 328350 282518 345922
rect 283052 423478 283108 423488
rect 283052 330958 283108 423422
rect 283052 330892 283108 330902
rect 284732 347172 284788 347182
rect 281898 328294 281994 328350
rect 282050 328294 282118 328350
rect 282174 328294 282242 328350
rect 282298 328294 282366 328350
rect 282422 328294 282518 328350
rect 281898 328226 282518 328294
rect 281898 328170 281994 328226
rect 282050 328170 282118 328226
rect 282174 328170 282242 328226
rect 282298 328170 282366 328226
rect 282422 328170 282518 328226
rect 281898 328102 282518 328170
rect 281898 328046 281994 328102
rect 282050 328046 282118 328102
rect 282174 328046 282242 328102
rect 282298 328046 282366 328102
rect 282422 328046 282518 328102
rect 281898 327978 282518 328046
rect 281898 327922 281994 327978
rect 282050 327922 282118 327978
rect 282174 327922 282242 327978
rect 282298 327922 282366 327978
rect 282422 327922 282518 327978
rect 278236 291778 278292 291788
rect 279692 313572 279748 313582
rect 277676 20132 277956 20188
rect 273868 14242 273924 14252
rect 270508 5954 270564 5964
rect 269388 5842 269444 5852
rect 267036 4274 267092 4284
rect 277900 4228 277956 20132
rect 279692 5124 279748 313516
rect 281372 312598 281428 312608
rect 281372 291956 281428 312542
rect 281372 291890 281428 291900
rect 281898 310350 282518 327922
rect 281898 310294 281994 310350
rect 282050 310294 282118 310350
rect 282174 310294 282242 310350
rect 282298 310294 282366 310350
rect 282422 310294 282518 310350
rect 281898 310226 282518 310294
rect 281898 310170 281994 310226
rect 282050 310170 282118 310226
rect 282174 310170 282242 310226
rect 282298 310170 282366 310226
rect 282422 310170 282518 310226
rect 281898 310102 282518 310170
rect 281898 310046 281994 310102
rect 282050 310046 282118 310102
rect 282174 310046 282242 310102
rect 282298 310046 282366 310102
rect 282422 310046 282518 310102
rect 281898 309978 282518 310046
rect 281898 309922 281994 309978
rect 282050 309922 282118 309978
rect 282174 309922 282242 309978
rect 282298 309922 282366 309978
rect 282422 309922 282518 309978
rect 281898 292350 282518 309922
rect 281898 292294 281994 292350
rect 282050 292294 282118 292350
rect 282174 292294 282242 292350
rect 282298 292294 282366 292350
rect 282422 292294 282518 292350
rect 281898 292226 282518 292294
rect 281898 292170 281994 292226
rect 282050 292170 282118 292226
rect 282174 292170 282242 292226
rect 282298 292170 282366 292226
rect 282422 292170 282518 292226
rect 281898 292102 282518 292170
rect 281898 292046 281994 292102
rect 282050 292046 282118 292102
rect 282174 292046 282242 292102
rect 282298 292046 282366 292102
rect 282422 292046 282518 292102
rect 281898 291978 282518 292046
rect 283052 321058 283108 321068
rect 283052 292068 283108 321002
rect 283052 292002 283108 292012
rect 281898 291922 281994 291978
rect 282050 291922 282118 291978
rect 282174 291922 282242 291978
rect 282298 291922 282366 291978
rect 282422 291922 282518 291978
rect 279692 5058 279748 5068
rect 281898 274350 282518 291922
rect 281898 274294 281994 274350
rect 282050 274294 282118 274350
rect 282174 274294 282242 274350
rect 282298 274294 282366 274350
rect 282422 274294 282518 274350
rect 281898 274226 282518 274294
rect 281898 274170 281994 274226
rect 282050 274170 282118 274226
rect 282174 274170 282242 274226
rect 282298 274170 282366 274226
rect 282422 274170 282518 274226
rect 281898 274102 282518 274170
rect 281898 274046 281994 274102
rect 282050 274046 282118 274102
rect 282174 274046 282242 274102
rect 282298 274046 282366 274102
rect 282422 274046 282518 274102
rect 281898 273978 282518 274046
rect 281898 273922 281994 273978
rect 282050 273922 282118 273978
rect 282174 273922 282242 273978
rect 282298 273922 282366 273978
rect 282422 273922 282518 273978
rect 281898 256350 282518 273922
rect 281898 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 282518 256350
rect 281898 256226 282518 256294
rect 281898 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 282518 256226
rect 281898 256102 282518 256170
rect 281898 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 282518 256102
rect 281898 255978 282518 256046
rect 281898 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 282518 255978
rect 281898 238350 282518 255922
rect 281898 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 282518 238350
rect 281898 238226 282518 238294
rect 281898 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 282518 238226
rect 281898 238102 282518 238170
rect 281898 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 282518 238102
rect 281898 237978 282518 238046
rect 281898 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 282518 237978
rect 281898 220350 282518 237922
rect 281898 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 282518 220350
rect 281898 220226 282518 220294
rect 281898 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 282518 220226
rect 281898 220102 282518 220170
rect 281898 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 282518 220102
rect 281898 219978 282518 220046
rect 281898 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 282518 219978
rect 281898 202350 282518 219922
rect 281898 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 282518 202350
rect 281898 202226 282518 202294
rect 281898 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 282518 202226
rect 281898 202102 282518 202170
rect 281898 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 282518 202102
rect 281898 201978 282518 202046
rect 281898 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 282518 201978
rect 281898 184350 282518 201922
rect 281898 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 282518 184350
rect 281898 184226 282518 184294
rect 281898 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 282518 184226
rect 281898 184102 282518 184170
rect 281898 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 282518 184102
rect 281898 183978 282518 184046
rect 281898 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 282518 183978
rect 281898 166350 282518 183922
rect 281898 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 282518 166350
rect 281898 166226 282518 166294
rect 281898 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 282518 166226
rect 281898 166102 282518 166170
rect 281898 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 282518 166102
rect 281898 165978 282518 166046
rect 281898 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 282518 165978
rect 281898 148350 282518 165922
rect 281898 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 282518 148350
rect 281898 148226 282518 148294
rect 281898 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 282518 148226
rect 281898 148102 282518 148170
rect 281898 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 282518 148102
rect 281898 147978 282518 148046
rect 281898 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 282518 147978
rect 281898 130350 282518 147922
rect 281898 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 282518 130350
rect 281898 130226 282518 130294
rect 281898 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 282518 130226
rect 281898 130102 282518 130170
rect 281898 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 282518 130102
rect 281898 129978 282518 130046
rect 281898 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 282518 129978
rect 281898 112350 282518 129922
rect 281898 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 282518 112350
rect 281898 112226 282518 112294
rect 281898 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 282518 112226
rect 281898 112102 282518 112170
rect 281898 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 282518 112102
rect 281898 111978 282518 112046
rect 281898 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 282518 111978
rect 281898 94350 282518 111922
rect 281898 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 282518 94350
rect 281898 94226 282518 94294
rect 281898 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 282518 94226
rect 281898 94102 282518 94170
rect 281898 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 282518 94102
rect 281898 93978 282518 94046
rect 281898 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 282518 93978
rect 281898 76350 282518 93922
rect 281898 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 282518 76350
rect 281898 76226 282518 76294
rect 281898 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 282518 76226
rect 281898 76102 282518 76170
rect 281898 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 282518 76102
rect 281898 75978 282518 76046
rect 281898 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 282518 75978
rect 281898 58350 282518 75922
rect 281898 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 282518 58350
rect 281898 58226 282518 58294
rect 281898 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 282518 58226
rect 281898 58102 282518 58170
rect 281898 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 282518 58102
rect 281898 57978 282518 58046
rect 281898 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 282518 57978
rect 281898 40350 282518 57922
rect 281898 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 282518 40350
rect 281898 40226 282518 40294
rect 281898 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 282518 40226
rect 281898 40102 282518 40170
rect 281898 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 282518 40102
rect 281898 39978 282518 40046
rect 281898 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 282518 39978
rect 281898 22350 282518 39922
rect 281898 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 282518 22350
rect 281898 22226 282518 22294
rect 281898 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 282518 22226
rect 281898 22102 282518 22170
rect 281898 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 282518 22102
rect 281898 21978 282518 22046
rect 281898 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 282518 21978
rect 277900 4162 277956 4172
rect 281898 4350 282518 21922
rect 284732 17668 284788 347116
rect 284844 206398 284900 429362
rect 284956 427364 285012 427374
rect 284956 345358 285012 427308
rect 284956 345292 285012 345302
rect 285618 424350 286238 441922
rect 288092 589798 288148 589808
rect 288092 437668 288148 589742
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 312618 562350 313238 579922
rect 312618 562294 312714 562350
rect 312770 562294 312838 562350
rect 312894 562294 312962 562350
rect 313018 562294 313086 562350
rect 313142 562294 313238 562350
rect 312618 562226 313238 562294
rect 312618 562170 312714 562226
rect 312770 562170 312838 562226
rect 312894 562170 312962 562226
rect 313018 562170 313086 562226
rect 313142 562170 313238 562226
rect 312618 562102 313238 562170
rect 312618 562046 312714 562102
rect 312770 562046 312838 562102
rect 312894 562046 312962 562102
rect 313018 562046 313086 562102
rect 313142 562046 313238 562102
rect 312618 561978 313238 562046
rect 312618 561922 312714 561978
rect 312770 561922 312838 561978
rect 312894 561922 312962 561978
rect 313018 561922 313086 561978
rect 313142 561922 313238 561978
rect 301084 550116 301140 550126
rect 300860 548884 300916 548894
rect 300748 546980 300804 546990
rect 300524 521780 300580 521796
rect 300524 521692 300580 521702
rect 300636 520324 300692 520356
rect 300636 520252 300692 520262
rect 300524 516898 300580 516908
rect 300524 516786 300580 516796
rect 300636 513658 300692 513668
rect 300636 513538 300692 513548
rect 300748 505876 300804 546924
rect 300860 511252 300916 548828
rect 300860 511186 300916 511196
rect 300972 547204 301028 547214
rect 300748 505810 300804 505820
rect 300972 503188 301028 547148
rect 301084 509068 301140 550060
rect 301756 550004 301812 550014
rect 301644 548548 301700 548558
rect 301532 547092 301588 547102
rect 301532 513658 301588 547036
rect 301644 516898 301700 548492
rect 301756 520318 301812 549948
rect 301868 549892 301924 549902
rect 301868 521758 301924 549836
rect 303436 548996 303492 549006
rect 301868 521692 301924 521702
rect 303212 548436 303268 548446
rect 301756 520252 301812 520262
rect 301644 516832 301700 516842
rect 301532 513592 301588 513602
rect 301084 509012 301588 509068
rect 300972 503122 301028 503132
rect 301532 502348 301588 509012
rect 301084 502292 301588 502348
rect 301084 497252 301140 502292
rect 301084 497186 301140 497196
rect 303212 472618 303268 548380
rect 303324 546868 303380 546878
rect 303324 488098 303380 546812
rect 303324 488032 303380 488042
rect 303436 479638 303492 548940
rect 312618 548142 313238 561922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 568350 316958 585922
rect 316338 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 316958 568350
rect 316338 568226 316958 568294
rect 316338 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 316958 568226
rect 316338 568102 316958 568170
rect 316338 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 316958 568102
rect 316338 567978 316958 568046
rect 316338 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 316958 567978
rect 316338 550350 316958 567922
rect 316338 550294 316434 550350
rect 316490 550294 316558 550350
rect 316614 550294 316682 550350
rect 316738 550294 316806 550350
rect 316862 550294 316958 550350
rect 316338 550226 316958 550294
rect 316338 550170 316434 550226
rect 316490 550170 316558 550226
rect 316614 550170 316682 550226
rect 316738 550170 316806 550226
rect 316862 550170 316958 550226
rect 316338 550102 316958 550170
rect 316338 550046 316434 550102
rect 316490 550046 316558 550102
rect 316614 550046 316682 550102
rect 316738 550046 316806 550102
rect 316862 550046 316958 550102
rect 316338 549978 316958 550046
rect 316338 549922 316434 549978
rect 316490 549922 316558 549978
rect 316614 549922 316682 549978
rect 316738 549922 316806 549978
rect 316862 549922 316958 549978
rect 316338 548142 316958 549922
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 343338 562350 343958 579922
rect 343338 562294 343434 562350
rect 343490 562294 343558 562350
rect 343614 562294 343682 562350
rect 343738 562294 343806 562350
rect 343862 562294 343958 562350
rect 343338 562226 343958 562294
rect 343338 562170 343434 562226
rect 343490 562170 343558 562226
rect 343614 562170 343682 562226
rect 343738 562170 343806 562226
rect 343862 562170 343958 562226
rect 343338 562102 343958 562170
rect 343338 562046 343434 562102
rect 343490 562046 343558 562102
rect 343614 562046 343682 562102
rect 343738 562046 343806 562102
rect 343862 562046 343958 562102
rect 343338 561978 343958 562046
rect 343338 561922 343434 561978
rect 343490 561922 343558 561978
rect 343614 561922 343682 561978
rect 343738 561922 343806 561978
rect 343862 561922 343958 561978
rect 323148 549444 323204 549454
rect 323148 548324 323204 549388
rect 323148 547204 323204 548268
rect 323148 547138 323204 547148
rect 328076 549444 328132 549454
rect 328076 546980 328132 549388
rect 333004 549444 333060 549454
rect 333004 549108 333060 549388
rect 333004 549042 333060 549052
rect 337932 549444 337988 549454
rect 337932 548436 337988 549388
rect 342860 549444 342916 549454
rect 342860 548996 342916 549388
rect 342860 548930 342916 548940
rect 337932 548370 337988 548380
rect 343338 548142 343958 561922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 568350 347678 585922
rect 347058 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 347678 568350
rect 347058 568226 347678 568294
rect 347058 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 347678 568226
rect 347058 568102 347678 568170
rect 347058 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 347678 568102
rect 347058 567978 347678 568046
rect 347058 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 347678 567978
rect 347058 550350 347678 567922
rect 347058 550294 347154 550350
rect 347210 550294 347278 550350
rect 347334 550294 347402 550350
rect 347458 550294 347526 550350
rect 347582 550294 347678 550350
rect 347058 550226 347678 550294
rect 347058 550170 347154 550226
rect 347210 550170 347278 550226
rect 347334 550170 347402 550226
rect 347458 550170 347526 550226
rect 347582 550170 347678 550226
rect 347058 550102 347678 550170
rect 347058 550046 347154 550102
rect 347210 550046 347278 550102
rect 347334 550046 347402 550102
rect 347458 550046 347526 550102
rect 347582 550046 347678 550102
rect 347058 549978 347678 550046
rect 347058 549922 347154 549978
rect 347210 549922 347278 549978
rect 347334 549922 347402 549978
rect 347458 549922 347526 549978
rect 347582 549922 347678 549978
rect 347058 548142 347678 549922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 374058 562350 374678 579922
rect 374058 562294 374154 562350
rect 374210 562294 374278 562350
rect 374334 562294 374402 562350
rect 374458 562294 374526 562350
rect 374582 562294 374678 562350
rect 374058 562226 374678 562294
rect 374058 562170 374154 562226
rect 374210 562170 374278 562226
rect 374334 562170 374402 562226
rect 374458 562170 374526 562226
rect 374582 562170 374678 562226
rect 374058 562102 374678 562170
rect 374058 562046 374154 562102
rect 374210 562046 374278 562102
rect 374334 562046 374402 562102
rect 374458 562046 374526 562102
rect 374582 562046 374678 562102
rect 374058 561978 374678 562046
rect 374058 561922 374154 561978
rect 374210 561922 374278 561978
rect 374334 561922 374402 561978
rect 374458 561922 374526 561978
rect 374582 561922 374678 561978
rect 362572 549556 362628 549566
rect 347788 549444 347844 549454
rect 328076 546914 328132 546924
rect 347788 546868 347844 549388
rect 352716 549444 352772 549454
rect 352716 548884 352772 549388
rect 352716 548818 352772 548828
rect 357644 549444 357700 549454
rect 357644 548436 357700 549388
rect 362572 548548 362628 549500
rect 362572 548482 362628 548492
rect 357644 547092 357700 548380
rect 374058 548142 374678 561922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 568350 378398 585922
rect 377778 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 378398 568350
rect 377778 568226 378398 568294
rect 377778 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 378398 568226
rect 377778 568102 378398 568170
rect 377778 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 378398 568102
rect 377778 567978 378398 568046
rect 377778 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 378398 567978
rect 377778 550350 378398 567922
rect 377778 550294 377874 550350
rect 377930 550294 377998 550350
rect 378054 550294 378122 550350
rect 378178 550294 378246 550350
rect 378302 550294 378398 550350
rect 377778 550226 378398 550294
rect 377778 550170 377874 550226
rect 377930 550170 377998 550226
rect 378054 550170 378122 550226
rect 378178 550170 378246 550226
rect 378302 550170 378398 550226
rect 377778 550102 378398 550170
rect 377778 550046 377874 550102
rect 377930 550046 377998 550102
rect 378054 550046 378122 550102
rect 378178 550046 378246 550102
rect 378302 550046 378398 550102
rect 377778 549978 378398 550046
rect 377778 549922 377874 549978
rect 377930 549922 377998 549978
rect 378054 549922 378122 549978
rect 378178 549922 378246 549978
rect 378302 549922 378398 549978
rect 377778 548142 378398 549922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 404778 562350 405398 579922
rect 404778 562294 404874 562350
rect 404930 562294 404998 562350
rect 405054 562294 405122 562350
rect 405178 562294 405246 562350
rect 405302 562294 405398 562350
rect 404778 562226 405398 562294
rect 404778 562170 404874 562226
rect 404930 562170 404998 562226
rect 405054 562170 405122 562226
rect 405178 562170 405246 562226
rect 405302 562170 405398 562226
rect 404778 562102 405398 562170
rect 404778 562046 404874 562102
rect 404930 562046 404998 562102
rect 405054 562046 405122 562102
rect 405178 562046 405246 562102
rect 405302 562046 405398 562102
rect 404778 561978 405398 562046
rect 404778 561922 404874 561978
rect 404930 561922 404998 561978
rect 405054 561922 405122 561978
rect 405178 561922 405246 561978
rect 405302 561922 405398 561978
rect 387212 549780 387268 549790
rect 386988 549220 387044 549230
rect 386988 548772 387044 549164
rect 386988 548706 387044 548716
rect 387212 548772 387268 549724
rect 392140 549444 392196 549454
rect 392140 549220 392196 549388
rect 392140 549154 392196 549164
rect 387212 548706 387268 548716
rect 404778 548142 405398 561922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 568350 409118 585922
rect 408498 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 409118 568350
rect 408498 568226 409118 568294
rect 408498 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 409118 568226
rect 408498 568102 409118 568170
rect 408498 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 409118 568102
rect 408498 567978 409118 568046
rect 408498 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 409118 567978
rect 408498 550350 409118 567922
rect 408498 550294 408594 550350
rect 408650 550294 408718 550350
rect 408774 550294 408842 550350
rect 408898 550294 408966 550350
rect 409022 550294 409118 550350
rect 408498 550226 409118 550294
rect 408498 550170 408594 550226
rect 408650 550170 408718 550226
rect 408774 550170 408842 550226
rect 408898 550170 408966 550226
rect 409022 550170 409118 550226
rect 408498 550102 409118 550170
rect 408498 550046 408594 550102
rect 408650 550046 408718 550102
rect 408774 550046 408842 550102
rect 408898 550046 408966 550102
rect 409022 550046 409118 550102
rect 408498 549978 409118 550046
rect 408498 549922 408594 549978
rect 408650 549922 408718 549978
rect 408774 549922 408842 549978
rect 408898 549922 408966 549978
rect 409022 549922 409118 549978
rect 408498 548142 409118 549922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 435498 562350 436118 579922
rect 435498 562294 435594 562350
rect 435650 562294 435718 562350
rect 435774 562294 435842 562350
rect 435898 562294 435966 562350
rect 436022 562294 436118 562350
rect 435498 562226 436118 562294
rect 435498 562170 435594 562226
rect 435650 562170 435718 562226
rect 435774 562170 435842 562226
rect 435898 562170 435966 562226
rect 436022 562170 436118 562226
rect 435498 562102 436118 562170
rect 435498 562046 435594 562102
rect 435650 562046 435718 562102
rect 435774 562046 435842 562102
rect 435898 562046 435966 562102
rect 436022 562046 436118 562102
rect 435498 561978 436118 562046
rect 435498 561922 435594 561978
rect 435650 561922 435718 561978
rect 435774 561922 435842 561978
rect 435898 561922 435966 561978
rect 436022 561922 436118 561978
rect 431676 549220 431732 549230
rect 431676 548772 431732 549164
rect 431676 548706 431732 548716
rect 435498 548142 436118 561922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 568350 439838 585922
rect 439218 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 439838 568350
rect 439218 568226 439838 568294
rect 439218 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 439838 568226
rect 439218 568102 439838 568170
rect 439218 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 439838 568102
rect 439218 567978 439838 568046
rect 439218 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 439838 567978
rect 439218 550350 439838 567922
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 466218 562350 466838 579922
rect 466218 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 466838 562350
rect 466218 562226 466838 562294
rect 466218 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 466838 562226
rect 466218 562102 466838 562170
rect 466218 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 466838 562102
rect 466218 561978 466838 562046
rect 466218 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 466838 561978
rect 459452 557938 459508 557948
rect 439218 550294 439314 550350
rect 439370 550294 439438 550350
rect 439494 550294 439562 550350
rect 439618 550294 439686 550350
rect 439742 550294 439838 550350
rect 439218 550226 439838 550294
rect 439218 550170 439314 550226
rect 439370 550170 439438 550226
rect 439494 550170 439562 550226
rect 439618 550170 439686 550226
rect 439742 550170 439838 550226
rect 439218 550102 439838 550170
rect 439218 550046 439314 550102
rect 439370 550046 439438 550102
rect 439494 550046 439562 550102
rect 439618 550046 439686 550102
rect 439742 550046 439838 550102
rect 439218 549978 439838 550046
rect 439218 549922 439314 549978
rect 439370 549922 439438 549978
rect 439494 549922 439562 549978
rect 439618 549922 439686 549978
rect 439742 549922 439838 549978
rect 439218 548142 439838 549922
rect 452732 551278 452788 551288
rect 446012 548772 446068 548782
rect 357644 547026 357700 547036
rect 347788 546802 347844 546812
rect 304448 544350 304768 544384
rect 304448 544294 304518 544350
rect 304574 544294 304642 544350
rect 304698 544294 304768 544350
rect 304448 544226 304768 544294
rect 304448 544170 304518 544226
rect 304574 544170 304642 544226
rect 304698 544170 304768 544226
rect 304448 544102 304768 544170
rect 304448 544046 304518 544102
rect 304574 544046 304642 544102
rect 304698 544046 304768 544102
rect 304448 543978 304768 544046
rect 304448 543922 304518 543978
rect 304574 543922 304642 543978
rect 304698 543922 304768 543978
rect 304448 543888 304768 543922
rect 335168 544350 335488 544384
rect 335168 544294 335238 544350
rect 335294 544294 335362 544350
rect 335418 544294 335488 544350
rect 335168 544226 335488 544294
rect 335168 544170 335238 544226
rect 335294 544170 335362 544226
rect 335418 544170 335488 544226
rect 335168 544102 335488 544170
rect 335168 544046 335238 544102
rect 335294 544046 335362 544102
rect 335418 544046 335488 544102
rect 335168 543978 335488 544046
rect 335168 543922 335238 543978
rect 335294 543922 335362 543978
rect 335418 543922 335488 543978
rect 335168 543888 335488 543922
rect 365888 544350 366208 544384
rect 365888 544294 365958 544350
rect 366014 544294 366082 544350
rect 366138 544294 366208 544350
rect 365888 544226 366208 544294
rect 365888 544170 365958 544226
rect 366014 544170 366082 544226
rect 366138 544170 366208 544226
rect 365888 544102 366208 544170
rect 365888 544046 365958 544102
rect 366014 544046 366082 544102
rect 366138 544046 366208 544102
rect 365888 543978 366208 544046
rect 365888 543922 365958 543978
rect 366014 543922 366082 543978
rect 366138 543922 366208 543978
rect 365888 543888 366208 543922
rect 396608 544350 396928 544384
rect 396608 544294 396678 544350
rect 396734 544294 396802 544350
rect 396858 544294 396928 544350
rect 396608 544226 396928 544294
rect 396608 544170 396678 544226
rect 396734 544170 396802 544226
rect 396858 544170 396928 544226
rect 396608 544102 396928 544170
rect 396608 544046 396678 544102
rect 396734 544046 396802 544102
rect 396858 544046 396928 544102
rect 396608 543978 396928 544046
rect 396608 543922 396678 543978
rect 396734 543922 396802 543978
rect 396858 543922 396928 543978
rect 396608 543888 396928 543922
rect 427328 544350 427648 544384
rect 427328 544294 427398 544350
rect 427454 544294 427522 544350
rect 427578 544294 427648 544350
rect 427328 544226 427648 544294
rect 427328 544170 427398 544226
rect 427454 544170 427522 544226
rect 427578 544170 427648 544226
rect 427328 544102 427648 544170
rect 427328 544046 427398 544102
rect 427454 544046 427522 544102
rect 427578 544046 427648 544102
rect 427328 543978 427648 544046
rect 427328 543922 427398 543978
rect 427454 543922 427522 543978
rect 427578 543922 427648 543978
rect 427328 543888 427648 543922
rect 319808 532350 320128 532384
rect 319808 532294 319878 532350
rect 319934 532294 320002 532350
rect 320058 532294 320128 532350
rect 319808 532226 320128 532294
rect 319808 532170 319878 532226
rect 319934 532170 320002 532226
rect 320058 532170 320128 532226
rect 319808 532102 320128 532170
rect 319808 532046 319878 532102
rect 319934 532046 320002 532102
rect 320058 532046 320128 532102
rect 319808 531978 320128 532046
rect 319808 531922 319878 531978
rect 319934 531922 320002 531978
rect 320058 531922 320128 531978
rect 319808 531888 320128 531922
rect 350528 532350 350848 532384
rect 350528 532294 350598 532350
rect 350654 532294 350722 532350
rect 350778 532294 350848 532350
rect 350528 532226 350848 532294
rect 350528 532170 350598 532226
rect 350654 532170 350722 532226
rect 350778 532170 350848 532226
rect 350528 532102 350848 532170
rect 350528 532046 350598 532102
rect 350654 532046 350722 532102
rect 350778 532046 350848 532102
rect 350528 531978 350848 532046
rect 350528 531922 350598 531978
rect 350654 531922 350722 531978
rect 350778 531922 350848 531978
rect 350528 531888 350848 531922
rect 381248 532350 381568 532384
rect 381248 532294 381318 532350
rect 381374 532294 381442 532350
rect 381498 532294 381568 532350
rect 381248 532226 381568 532294
rect 381248 532170 381318 532226
rect 381374 532170 381442 532226
rect 381498 532170 381568 532226
rect 381248 532102 381568 532170
rect 381248 532046 381318 532102
rect 381374 532046 381442 532102
rect 381498 532046 381568 532102
rect 381248 531978 381568 532046
rect 381248 531922 381318 531978
rect 381374 531922 381442 531978
rect 381498 531922 381568 531978
rect 381248 531888 381568 531922
rect 411968 532350 412288 532384
rect 411968 532294 412038 532350
rect 412094 532294 412162 532350
rect 412218 532294 412288 532350
rect 411968 532226 412288 532294
rect 411968 532170 412038 532226
rect 412094 532170 412162 532226
rect 412218 532170 412288 532226
rect 411968 532102 412288 532170
rect 411968 532046 412038 532102
rect 412094 532046 412162 532102
rect 412218 532046 412288 532102
rect 411968 531978 412288 532046
rect 411968 531922 412038 531978
rect 412094 531922 412162 531978
rect 412218 531922 412288 531978
rect 411968 531888 412288 531922
rect 442688 532350 443008 532384
rect 442688 532294 442758 532350
rect 442814 532294 442882 532350
rect 442938 532294 443008 532350
rect 442688 532226 443008 532294
rect 442688 532170 442758 532226
rect 442814 532170 442882 532226
rect 442938 532170 443008 532226
rect 442688 532102 443008 532170
rect 442688 532046 442758 532102
rect 442814 532046 442882 532102
rect 442938 532046 443008 532102
rect 442688 531978 443008 532046
rect 442688 531922 442758 531978
rect 442814 531922 442882 531978
rect 442938 531922 443008 531978
rect 442688 531888 443008 531922
rect 304448 526350 304768 526384
rect 304448 526294 304518 526350
rect 304574 526294 304642 526350
rect 304698 526294 304768 526350
rect 304448 526226 304768 526294
rect 304448 526170 304518 526226
rect 304574 526170 304642 526226
rect 304698 526170 304768 526226
rect 304448 526102 304768 526170
rect 304448 526046 304518 526102
rect 304574 526046 304642 526102
rect 304698 526046 304768 526102
rect 304448 525978 304768 526046
rect 304448 525922 304518 525978
rect 304574 525922 304642 525978
rect 304698 525922 304768 525978
rect 304448 525888 304768 525922
rect 335168 526350 335488 526384
rect 335168 526294 335238 526350
rect 335294 526294 335362 526350
rect 335418 526294 335488 526350
rect 335168 526226 335488 526294
rect 335168 526170 335238 526226
rect 335294 526170 335362 526226
rect 335418 526170 335488 526226
rect 335168 526102 335488 526170
rect 335168 526046 335238 526102
rect 335294 526046 335362 526102
rect 335418 526046 335488 526102
rect 335168 525978 335488 526046
rect 335168 525922 335238 525978
rect 335294 525922 335362 525978
rect 335418 525922 335488 525978
rect 335168 525888 335488 525922
rect 365888 526350 366208 526384
rect 365888 526294 365958 526350
rect 366014 526294 366082 526350
rect 366138 526294 366208 526350
rect 365888 526226 366208 526294
rect 365888 526170 365958 526226
rect 366014 526170 366082 526226
rect 366138 526170 366208 526226
rect 365888 526102 366208 526170
rect 365888 526046 365958 526102
rect 366014 526046 366082 526102
rect 366138 526046 366208 526102
rect 365888 525978 366208 526046
rect 365888 525922 365958 525978
rect 366014 525922 366082 525978
rect 366138 525922 366208 525978
rect 365888 525888 366208 525922
rect 396608 526350 396928 526384
rect 396608 526294 396678 526350
rect 396734 526294 396802 526350
rect 396858 526294 396928 526350
rect 396608 526226 396928 526294
rect 396608 526170 396678 526226
rect 396734 526170 396802 526226
rect 396858 526170 396928 526226
rect 396608 526102 396928 526170
rect 396608 526046 396678 526102
rect 396734 526046 396802 526102
rect 396858 526046 396928 526102
rect 396608 525978 396928 526046
rect 396608 525922 396678 525978
rect 396734 525922 396802 525978
rect 396858 525922 396928 525978
rect 396608 525888 396928 525922
rect 427328 526350 427648 526384
rect 427328 526294 427398 526350
rect 427454 526294 427522 526350
rect 427578 526294 427648 526350
rect 427328 526226 427648 526294
rect 427328 526170 427398 526226
rect 427454 526170 427522 526226
rect 427578 526170 427648 526226
rect 427328 526102 427648 526170
rect 427328 526046 427398 526102
rect 427454 526046 427522 526102
rect 427578 526046 427648 526102
rect 427328 525978 427648 526046
rect 427328 525922 427398 525978
rect 427454 525922 427522 525978
rect 427578 525922 427648 525978
rect 427328 525888 427648 525922
rect 319808 514350 320128 514384
rect 319808 514294 319878 514350
rect 319934 514294 320002 514350
rect 320058 514294 320128 514350
rect 319808 514226 320128 514294
rect 319808 514170 319878 514226
rect 319934 514170 320002 514226
rect 320058 514170 320128 514226
rect 319808 514102 320128 514170
rect 319808 514046 319878 514102
rect 319934 514046 320002 514102
rect 320058 514046 320128 514102
rect 319808 513978 320128 514046
rect 319808 513922 319878 513978
rect 319934 513922 320002 513978
rect 320058 513922 320128 513978
rect 319808 513888 320128 513922
rect 350528 514350 350848 514384
rect 350528 514294 350598 514350
rect 350654 514294 350722 514350
rect 350778 514294 350848 514350
rect 350528 514226 350848 514294
rect 350528 514170 350598 514226
rect 350654 514170 350722 514226
rect 350778 514170 350848 514226
rect 350528 514102 350848 514170
rect 350528 514046 350598 514102
rect 350654 514046 350722 514102
rect 350778 514046 350848 514102
rect 350528 513978 350848 514046
rect 350528 513922 350598 513978
rect 350654 513922 350722 513978
rect 350778 513922 350848 513978
rect 350528 513888 350848 513922
rect 381248 514350 381568 514384
rect 381248 514294 381318 514350
rect 381374 514294 381442 514350
rect 381498 514294 381568 514350
rect 381248 514226 381568 514294
rect 381248 514170 381318 514226
rect 381374 514170 381442 514226
rect 381498 514170 381568 514226
rect 381248 514102 381568 514170
rect 381248 514046 381318 514102
rect 381374 514046 381442 514102
rect 381498 514046 381568 514102
rect 381248 513978 381568 514046
rect 381248 513922 381318 513978
rect 381374 513922 381442 513978
rect 381498 513922 381568 513978
rect 381248 513888 381568 513922
rect 411968 514350 412288 514384
rect 411968 514294 412038 514350
rect 412094 514294 412162 514350
rect 412218 514294 412288 514350
rect 411968 514226 412288 514294
rect 411968 514170 412038 514226
rect 412094 514170 412162 514226
rect 412218 514170 412288 514226
rect 411968 514102 412288 514170
rect 411968 514046 412038 514102
rect 412094 514046 412162 514102
rect 412218 514046 412288 514102
rect 411968 513978 412288 514046
rect 411968 513922 412038 513978
rect 412094 513922 412162 513978
rect 412218 513922 412288 513978
rect 411968 513888 412288 513922
rect 442688 514350 443008 514384
rect 442688 514294 442758 514350
rect 442814 514294 442882 514350
rect 442938 514294 443008 514350
rect 442688 514226 443008 514294
rect 442688 514170 442758 514226
rect 442814 514170 442882 514226
rect 442938 514170 443008 514226
rect 442688 514102 443008 514170
rect 442688 514046 442758 514102
rect 442814 514046 442882 514102
rect 442938 514046 443008 514102
rect 442688 513978 443008 514046
rect 442688 513922 442758 513978
rect 442814 513922 442882 513978
rect 442938 513922 443008 513978
rect 442688 513888 443008 513922
rect 304448 508350 304768 508384
rect 304448 508294 304518 508350
rect 304574 508294 304642 508350
rect 304698 508294 304768 508350
rect 304448 508226 304768 508294
rect 304448 508170 304518 508226
rect 304574 508170 304642 508226
rect 304698 508170 304768 508226
rect 304448 508102 304768 508170
rect 304448 508046 304518 508102
rect 304574 508046 304642 508102
rect 304698 508046 304768 508102
rect 304448 507978 304768 508046
rect 304448 507922 304518 507978
rect 304574 507922 304642 507978
rect 304698 507922 304768 507978
rect 304448 507888 304768 507922
rect 335168 508350 335488 508384
rect 335168 508294 335238 508350
rect 335294 508294 335362 508350
rect 335418 508294 335488 508350
rect 335168 508226 335488 508294
rect 335168 508170 335238 508226
rect 335294 508170 335362 508226
rect 335418 508170 335488 508226
rect 335168 508102 335488 508170
rect 335168 508046 335238 508102
rect 335294 508046 335362 508102
rect 335418 508046 335488 508102
rect 335168 507978 335488 508046
rect 335168 507922 335238 507978
rect 335294 507922 335362 507978
rect 335418 507922 335488 507978
rect 335168 507888 335488 507922
rect 365888 508350 366208 508384
rect 365888 508294 365958 508350
rect 366014 508294 366082 508350
rect 366138 508294 366208 508350
rect 365888 508226 366208 508294
rect 365888 508170 365958 508226
rect 366014 508170 366082 508226
rect 366138 508170 366208 508226
rect 365888 508102 366208 508170
rect 365888 508046 365958 508102
rect 366014 508046 366082 508102
rect 366138 508046 366208 508102
rect 365888 507978 366208 508046
rect 365888 507922 365958 507978
rect 366014 507922 366082 507978
rect 366138 507922 366208 507978
rect 365888 507888 366208 507922
rect 396608 508350 396928 508384
rect 396608 508294 396678 508350
rect 396734 508294 396802 508350
rect 396858 508294 396928 508350
rect 396608 508226 396928 508294
rect 396608 508170 396678 508226
rect 396734 508170 396802 508226
rect 396858 508170 396928 508226
rect 396608 508102 396928 508170
rect 396608 508046 396678 508102
rect 396734 508046 396802 508102
rect 396858 508046 396928 508102
rect 396608 507978 396928 508046
rect 396608 507922 396678 507978
rect 396734 507922 396802 507978
rect 396858 507922 396928 507978
rect 396608 507888 396928 507922
rect 427328 508350 427648 508384
rect 427328 508294 427398 508350
rect 427454 508294 427522 508350
rect 427578 508294 427648 508350
rect 427328 508226 427648 508294
rect 427328 508170 427398 508226
rect 427454 508170 427522 508226
rect 427578 508170 427648 508226
rect 427328 508102 427648 508170
rect 427328 508046 427398 508102
rect 427454 508046 427522 508102
rect 427578 508046 427648 508102
rect 427328 507978 427648 508046
rect 427328 507922 427398 507978
rect 427454 507922 427522 507978
rect 427578 507922 427648 507978
rect 427328 507888 427648 507922
rect 446012 499798 446068 548716
rect 446012 499732 446068 499742
rect 319808 496350 320128 496384
rect 319808 496294 319878 496350
rect 319934 496294 320002 496350
rect 320058 496294 320128 496350
rect 319808 496226 320128 496294
rect 319808 496170 319878 496226
rect 319934 496170 320002 496226
rect 320058 496170 320128 496226
rect 319808 496102 320128 496170
rect 319808 496046 319878 496102
rect 319934 496046 320002 496102
rect 320058 496046 320128 496102
rect 319808 495978 320128 496046
rect 319808 495922 319878 495978
rect 319934 495922 320002 495978
rect 320058 495922 320128 495978
rect 319808 495888 320128 495922
rect 350528 496350 350848 496384
rect 350528 496294 350598 496350
rect 350654 496294 350722 496350
rect 350778 496294 350848 496350
rect 350528 496226 350848 496294
rect 350528 496170 350598 496226
rect 350654 496170 350722 496226
rect 350778 496170 350848 496226
rect 350528 496102 350848 496170
rect 350528 496046 350598 496102
rect 350654 496046 350722 496102
rect 350778 496046 350848 496102
rect 350528 495978 350848 496046
rect 350528 495922 350598 495978
rect 350654 495922 350722 495978
rect 350778 495922 350848 495978
rect 350528 495888 350848 495922
rect 381248 496350 381568 496384
rect 381248 496294 381318 496350
rect 381374 496294 381442 496350
rect 381498 496294 381568 496350
rect 381248 496226 381568 496294
rect 381248 496170 381318 496226
rect 381374 496170 381442 496226
rect 381498 496170 381568 496226
rect 381248 496102 381568 496170
rect 381248 496046 381318 496102
rect 381374 496046 381442 496102
rect 381498 496046 381568 496102
rect 381248 495978 381568 496046
rect 381248 495922 381318 495978
rect 381374 495922 381442 495978
rect 381498 495922 381568 495978
rect 381248 495888 381568 495922
rect 411968 496350 412288 496384
rect 411968 496294 412038 496350
rect 412094 496294 412162 496350
rect 412218 496294 412288 496350
rect 411968 496226 412288 496294
rect 411968 496170 412038 496226
rect 412094 496170 412162 496226
rect 412218 496170 412288 496226
rect 411968 496102 412288 496170
rect 411968 496046 412038 496102
rect 412094 496046 412162 496102
rect 412218 496046 412288 496102
rect 411968 495978 412288 496046
rect 411968 495922 412038 495978
rect 412094 495922 412162 495978
rect 412218 495922 412288 495978
rect 411968 495888 412288 495922
rect 442688 496350 443008 496384
rect 442688 496294 442758 496350
rect 442814 496294 442882 496350
rect 442938 496294 443008 496350
rect 442688 496226 443008 496294
rect 442688 496170 442758 496226
rect 442814 496170 442882 496226
rect 442938 496170 443008 496226
rect 442688 496102 443008 496170
rect 442688 496046 442758 496102
rect 442814 496046 442882 496102
rect 442938 496046 443008 496102
rect 442688 495978 443008 496046
rect 442688 495922 442758 495978
rect 442814 495922 442882 495978
rect 442938 495922 443008 495978
rect 442688 495888 443008 495922
rect 304448 490350 304768 490384
rect 304448 490294 304518 490350
rect 304574 490294 304642 490350
rect 304698 490294 304768 490350
rect 304448 490226 304768 490294
rect 304448 490170 304518 490226
rect 304574 490170 304642 490226
rect 304698 490170 304768 490226
rect 304448 490102 304768 490170
rect 304448 490046 304518 490102
rect 304574 490046 304642 490102
rect 304698 490046 304768 490102
rect 304448 489978 304768 490046
rect 304448 489922 304518 489978
rect 304574 489922 304642 489978
rect 304698 489922 304768 489978
rect 304448 489888 304768 489922
rect 335168 490350 335488 490384
rect 335168 490294 335238 490350
rect 335294 490294 335362 490350
rect 335418 490294 335488 490350
rect 335168 490226 335488 490294
rect 335168 490170 335238 490226
rect 335294 490170 335362 490226
rect 335418 490170 335488 490226
rect 335168 490102 335488 490170
rect 335168 490046 335238 490102
rect 335294 490046 335362 490102
rect 335418 490046 335488 490102
rect 335168 489978 335488 490046
rect 335168 489922 335238 489978
rect 335294 489922 335362 489978
rect 335418 489922 335488 489978
rect 335168 489888 335488 489922
rect 365888 490350 366208 490384
rect 365888 490294 365958 490350
rect 366014 490294 366082 490350
rect 366138 490294 366208 490350
rect 365888 490226 366208 490294
rect 365888 490170 365958 490226
rect 366014 490170 366082 490226
rect 366138 490170 366208 490226
rect 365888 490102 366208 490170
rect 365888 490046 365958 490102
rect 366014 490046 366082 490102
rect 366138 490046 366208 490102
rect 365888 489978 366208 490046
rect 365888 489922 365958 489978
rect 366014 489922 366082 489978
rect 366138 489922 366208 489978
rect 365888 489888 366208 489922
rect 396608 490350 396928 490384
rect 396608 490294 396678 490350
rect 396734 490294 396802 490350
rect 396858 490294 396928 490350
rect 396608 490226 396928 490294
rect 396608 490170 396678 490226
rect 396734 490170 396802 490226
rect 396858 490170 396928 490226
rect 396608 490102 396928 490170
rect 396608 490046 396678 490102
rect 396734 490046 396802 490102
rect 396858 490046 396928 490102
rect 396608 489978 396928 490046
rect 396608 489922 396678 489978
rect 396734 489922 396802 489978
rect 396858 489922 396928 489978
rect 396608 489888 396928 489922
rect 427328 490350 427648 490384
rect 427328 490294 427398 490350
rect 427454 490294 427522 490350
rect 427578 490294 427648 490350
rect 427328 490226 427648 490294
rect 427328 490170 427398 490226
rect 427454 490170 427522 490226
rect 427578 490170 427648 490226
rect 427328 490102 427648 490170
rect 427328 490046 427398 490102
rect 427454 490046 427522 490102
rect 427578 490046 427648 490102
rect 427328 489978 427648 490046
rect 427328 489922 427398 489978
rect 427454 489922 427522 489978
rect 427578 489922 427648 489978
rect 427328 489888 427648 489922
rect 303436 479572 303492 479582
rect 319808 478350 320128 478384
rect 319808 478294 319878 478350
rect 319934 478294 320002 478350
rect 320058 478294 320128 478350
rect 319808 478226 320128 478294
rect 319808 478170 319878 478226
rect 319934 478170 320002 478226
rect 320058 478170 320128 478226
rect 319808 478102 320128 478170
rect 319808 478046 319878 478102
rect 319934 478046 320002 478102
rect 320058 478046 320128 478102
rect 319808 477978 320128 478046
rect 319808 477922 319878 477978
rect 319934 477922 320002 477978
rect 320058 477922 320128 477978
rect 319808 477888 320128 477922
rect 350528 478350 350848 478384
rect 350528 478294 350598 478350
rect 350654 478294 350722 478350
rect 350778 478294 350848 478350
rect 350528 478226 350848 478294
rect 350528 478170 350598 478226
rect 350654 478170 350722 478226
rect 350778 478170 350848 478226
rect 350528 478102 350848 478170
rect 350528 478046 350598 478102
rect 350654 478046 350722 478102
rect 350778 478046 350848 478102
rect 350528 477978 350848 478046
rect 350528 477922 350598 477978
rect 350654 477922 350722 477978
rect 350778 477922 350848 477978
rect 350528 477888 350848 477922
rect 381248 478350 381568 478384
rect 381248 478294 381318 478350
rect 381374 478294 381442 478350
rect 381498 478294 381568 478350
rect 381248 478226 381568 478294
rect 381248 478170 381318 478226
rect 381374 478170 381442 478226
rect 381498 478170 381568 478226
rect 381248 478102 381568 478170
rect 381248 478046 381318 478102
rect 381374 478046 381442 478102
rect 381498 478046 381568 478102
rect 381248 477978 381568 478046
rect 381248 477922 381318 477978
rect 381374 477922 381442 477978
rect 381498 477922 381568 477978
rect 381248 477888 381568 477922
rect 411968 478350 412288 478384
rect 411968 478294 412038 478350
rect 412094 478294 412162 478350
rect 412218 478294 412288 478350
rect 411968 478226 412288 478294
rect 411968 478170 412038 478226
rect 412094 478170 412162 478226
rect 412218 478170 412288 478226
rect 411968 478102 412288 478170
rect 411968 478046 412038 478102
rect 412094 478046 412162 478102
rect 412218 478046 412288 478102
rect 411968 477978 412288 478046
rect 411968 477922 412038 477978
rect 412094 477922 412162 477978
rect 412218 477922 412288 477978
rect 411968 477888 412288 477922
rect 442688 478350 443008 478384
rect 442688 478294 442758 478350
rect 442814 478294 442882 478350
rect 442938 478294 443008 478350
rect 442688 478226 443008 478294
rect 442688 478170 442758 478226
rect 442814 478170 442882 478226
rect 442938 478170 443008 478226
rect 442688 478102 443008 478170
rect 442688 478046 442758 478102
rect 442814 478046 442882 478102
rect 442938 478046 443008 478102
rect 442688 477978 443008 478046
rect 442688 477922 442758 477978
rect 442814 477922 442882 477978
rect 442938 477922 443008 477978
rect 442688 477888 443008 477922
rect 288092 437602 288148 437612
rect 293132 452788 293188 452798
rect 288204 431938 288260 431948
rect 285618 424294 285714 424350
rect 285770 424294 285838 424350
rect 285894 424294 285962 424350
rect 286018 424294 286086 424350
rect 286142 424294 286238 424350
rect 285618 424226 286238 424294
rect 285618 424170 285714 424226
rect 285770 424170 285838 424226
rect 285894 424170 285962 424226
rect 286018 424170 286086 424226
rect 286142 424170 286238 424226
rect 285618 424102 286238 424170
rect 285618 424046 285714 424102
rect 285770 424046 285838 424102
rect 285894 424046 285962 424102
rect 286018 424046 286086 424102
rect 286142 424046 286238 424102
rect 285618 423978 286238 424046
rect 285618 423922 285714 423978
rect 285770 423922 285838 423978
rect 285894 423922 285962 423978
rect 286018 423922 286086 423978
rect 286142 423922 286238 423978
rect 285618 406350 286238 423922
rect 285618 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 286238 406350
rect 285618 406226 286238 406294
rect 285618 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 286238 406226
rect 285618 406102 286238 406170
rect 285618 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 286238 406102
rect 285618 405978 286238 406046
rect 285618 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 286238 405978
rect 285618 388350 286238 405922
rect 285618 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 286238 388350
rect 285618 388226 286238 388294
rect 285618 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 286238 388226
rect 285618 388102 286238 388170
rect 285618 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 286238 388102
rect 285618 387978 286238 388046
rect 285618 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 286238 387978
rect 285618 370350 286238 387922
rect 285618 370294 285714 370350
rect 285770 370294 285838 370350
rect 285894 370294 285962 370350
rect 286018 370294 286086 370350
rect 286142 370294 286238 370350
rect 285618 370226 286238 370294
rect 285618 370170 285714 370226
rect 285770 370170 285838 370226
rect 285894 370170 285962 370226
rect 286018 370170 286086 370226
rect 286142 370170 286238 370226
rect 285618 370102 286238 370170
rect 285618 370046 285714 370102
rect 285770 370046 285838 370102
rect 285894 370046 285962 370102
rect 286018 370046 286086 370102
rect 286142 370046 286238 370102
rect 285618 369978 286238 370046
rect 285618 369922 285714 369978
rect 285770 369922 285838 369978
rect 285894 369922 285962 369978
rect 286018 369922 286086 369978
rect 286142 369922 286238 369978
rect 285618 352350 286238 369922
rect 285618 352294 285714 352350
rect 285770 352294 285838 352350
rect 285894 352294 285962 352350
rect 286018 352294 286086 352350
rect 286142 352294 286238 352350
rect 285618 352226 286238 352294
rect 285618 352170 285714 352226
rect 285770 352170 285838 352226
rect 285894 352170 285962 352226
rect 286018 352170 286086 352226
rect 286142 352170 286238 352226
rect 285618 352102 286238 352170
rect 285618 352046 285714 352102
rect 285770 352046 285838 352102
rect 285894 352046 285962 352102
rect 286018 352046 286086 352102
rect 286142 352046 286238 352102
rect 285618 351978 286238 352046
rect 285618 351922 285714 351978
rect 285770 351922 285838 351978
rect 285894 351922 285962 351978
rect 286018 351922 286086 351978
rect 286142 351922 286238 351978
rect 284844 206332 284900 206342
rect 285618 334350 286238 351922
rect 288092 430724 288148 430734
rect 288092 339238 288148 430668
rect 288092 339172 288148 339182
rect 285618 334294 285714 334350
rect 285770 334294 285838 334350
rect 285894 334294 285962 334350
rect 286018 334294 286086 334350
rect 286142 334294 286238 334350
rect 285618 334226 286238 334294
rect 285618 334170 285714 334226
rect 285770 334170 285838 334226
rect 285894 334170 285962 334226
rect 286018 334170 286086 334226
rect 286142 334170 286238 334226
rect 285618 334102 286238 334170
rect 285618 334046 285714 334102
rect 285770 334046 285838 334102
rect 285894 334046 285962 334102
rect 286018 334046 286086 334102
rect 286142 334046 286238 334102
rect 285618 333978 286238 334046
rect 285618 333922 285714 333978
rect 285770 333922 285838 333978
rect 285894 333922 285962 333978
rect 286018 333922 286086 333978
rect 286142 333922 286238 333978
rect 285618 316350 286238 333922
rect 285618 316294 285714 316350
rect 285770 316294 285838 316350
rect 285894 316294 285962 316350
rect 286018 316294 286086 316350
rect 286142 316294 286238 316350
rect 285618 316226 286238 316294
rect 285618 316170 285714 316226
rect 285770 316170 285838 316226
rect 285894 316170 285962 316226
rect 286018 316170 286086 316226
rect 286142 316170 286238 316226
rect 285618 316102 286238 316170
rect 285618 316046 285714 316102
rect 285770 316046 285838 316102
rect 285894 316046 285962 316102
rect 286018 316046 286086 316102
rect 286142 316046 286238 316102
rect 285618 315978 286238 316046
rect 285618 315922 285714 315978
rect 285770 315922 285838 315978
rect 285894 315922 285962 315978
rect 286018 315922 286086 315978
rect 286142 315922 286238 315978
rect 285618 298350 286238 315922
rect 285618 298294 285714 298350
rect 285770 298294 285838 298350
rect 285894 298294 285962 298350
rect 286018 298294 286086 298350
rect 286142 298294 286238 298350
rect 285618 298226 286238 298294
rect 285618 298170 285714 298226
rect 285770 298170 285838 298226
rect 285894 298170 285962 298226
rect 286018 298170 286086 298226
rect 286142 298170 286238 298226
rect 285618 298102 286238 298170
rect 285618 298046 285714 298102
rect 285770 298046 285838 298102
rect 285894 298046 285962 298102
rect 286018 298046 286086 298102
rect 286142 298046 286238 298102
rect 285618 297978 286238 298046
rect 285618 297922 285714 297978
rect 285770 297922 285838 297978
rect 285894 297922 285962 297978
rect 286018 297922 286086 297978
rect 286142 297922 286238 297978
rect 285618 280350 286238 297922
rect 285618 280294 285714 280350
rect 285770 280294 285838 280350
rect 285894 280294 285962 280350
rect 286018 280294 286086 280350
rect 286142 280294 286238 280350
rect 285618 280226 286238 280294
rect 285618 280170 285714 280226
rect 285770 280170 285838 280226
rect 285894 280170 285962 280226
rect 286018 280170 286086 280226
rect 286142 280170 286238 280226
rect 285618 280102 286238 280170
rect 285618 280046 285714 280102
rect 285770 280046 285838 280102
rect 285894 280046 285962 280102
rect 286018 280046 286086 280102
rect 286142 280046 286238 280102
rect 285618 279978 286238 280046
rect 285618 279922 285714 279978
rect 285770 279922 285838 279978
rect 285894 279922 285962 279978
rect 286018 279922 286086 279978
rect 286142 279922 286238 279978
rect 285618 262350 286238 279922
rect 285618 262294 285714 262350
rect 285770 262294 285838 262350
rect 285894 262294 285962 262350
rect 286018 262294 286086 262350
rect 286142 262294 286238 262350
rect 285618 262226 286238 262294
rect 285618 262170 285714 262226
rect 285770 262170 285838 262226
rect 285894 262170 285962 262226
rect 286018 262170 286086 262226
rect 286142 262170 286238 262226
rect 285618 262102 286238 262170
rect 285618 262046 285714 262102
rect 285770 262046 285838 262102
rect 285894 262046 285962 262102
rect 286018 262046 286086 262102
rect 286142 262046 286238 262102
rect 285618 261978 286238 262046
rect 285618 261922 285714 261978
rect 285770 261922 285838 261978
rect 285894 261922 285962 261978
rect 286018 261922 286086 261978
rect 286142 261922 286238 261978
rect 285618 244350 286238 261922
rect 285618 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 286238 244350
rect 285618 244226 286238 244294
rect 285618 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 286238 244226
rect 285618 244102 286238 244170
rect 285618 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 286238 244102
rect 285618 243978 286238 244046
rect 285618 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 286238 243978
rect 285618 226350 286238 243922
rect 285618 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 286238 226350
rect 285618 226226 286238 226294
rect 285618 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 286238 226226
rect 285618 226102 286238 226170
rect 285618 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 286238 226102
rect 285618 225978 286238 226046
rect 285618 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 286238 225978
rect 285618 208350 286238 225922
rect 285618 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 286238 208350
rect 285618 208226 286238 208294
rect 285618 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 286238 208226
rect 285618 208102 286238 208170
rect 285618 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 286238 208102
rect 285618 207978 286238 208046
rect 285618 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 286238 207978
rect 284732 17602 284788 17612
rect 285618 190350 286238 207922
rect 285618 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 286238 190350
rect 285618 190226 286238 190294
rect 285618 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 286238 190226
rect 285618 190102 286238 190170
rect 285618 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 286238 190102
rect 285618 189978 286238 190046
rect 285618 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 286238 189978
rect 285618 172350 286238 189922
rect 285618 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 286238 172350
rect 285618 172226 286238 172294
rect 285618 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 286238 172226
rect 285618 172102 286238 172170
rect 285618 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 286238 172102
rect 285618 171978 286238 172046
rect 285618 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 286238 171978
rect 285618 154350 286238 171922
rect 285618 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 286238 154350
rect 285618 154226 286238 154294
rect 285618 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 286238 154226
rect 285618 154102 286238 154170
rect 285618 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 286238 154102
rect 285618 153978 286238 154046
rect 285618 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 286238 153978
rect 285618 136350 286238 153922
rect 285618 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 286238 136350
rect 285618 136226 286238 136294
rect 285618 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 286238 136226
rect 285618 136102 286238 136170
rect 285618 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 286238 136102
rect 285618 135978 286238 136046
rect 285618 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 286238 135978
rect 285618 118350 286238 135922
rect 285618 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 286238 118350
rect 285618 118226 286238 118294
rect 285618 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 286238 118226
rect 285618 118102 286238 118170
rect 285618 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 286238 118102
rect 285618 117978 286238 118046
rect 285618 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 286238 117978
rect 285618 100350 286238 117922
rect 285618 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 286238 100350
rect 285618 100226 286238 100294
rect 285618 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 286238 100226
rect 285618 100102 286238 100170
rect 285618 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 286238 100102
rect 285618 99978 286238 100046
rect 285618 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 286238 99978
rect 285618 82350 286238 99922
rect 285618 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 286238 82350
rect 285618 82226 286238 82294
rect 285618 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 286238 82226
rect 285618 82102 286238 82170
rect 285618 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 286238 82102
rect 285618 81978 286238 82046
rect 285618 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 286238 81978
rect 285618 64350 286238 81922
rect 285618 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 286238 64350
rect 285618 64226 286238 64294
rect 285618 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 286238 64226
rect 285618 64102 286238 64170
rect 285618 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 286238 64102
rect 285618 63978 286238 64046
rect 285618 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 286238 63978
rect 285618 46350 286238 63922
rect 285618 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 286238 46350
rect 285618 46226 286238 46294
rect 285618 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 286238 46226
rect 285618 46102 286238 46170
rect 285618 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 286238 46102
rect 285618 45978 286238 46046
rect 285618 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 286238 45978
rect 285618 28350 286238 45922
rect 285618 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 286238 28350
rect 285618 28226 286238 28294
rect 285618 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 286238 28226
rect 285618 28102 286238 28170
rect 285618 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 286238 28102
rect 285618 27978 286238 28046
rect 285618 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 286238 27978
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 285618 10350 286238 27922
rect 285618 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 286238 10350
rect 285618 10226 286238 10294
rect 285618 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 286238 10226
rect 285618 10102 286238 10170
rect 285618 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 286238 10102
rect 285618 9978 286238 10046
rect 285618 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 286238 9978
rect 285618 -1120 286238 9922
rect 288092 314916 288148 314926
rect 288092 5124 288148 314860
rect 288204 268100 288260 431882
rect 291564 429492 291620 429502
rect 289884 429268 289940 429278
rect 289772 427078 289828 427088
rect 289772 345538 289828 427022
rect 289884 377938 289940 429212
rect 289884 377872 289940 377882
rect 289772 345472 289828 345482
rect 291452 345828 291508 345838
rect 288316 326098 288372 326108
rect 288316 292740 288372 326042
rect 289884 317818 289940 317828
rect 288316 292674 288372 292684
rect 289772 316260 289828 316270
rect 288204 268034 288260 268044
rect 289772 6020 289828 316204
rect 289884 292180 289940 317762
rect 289884 292114 289940 292124
rect 291452 15988 291508 345772
rect 291564 285238 291620 429436
rect 293132 377758 293188 452732
rect 298396 436212 298452 436222
rect 296604 430858 296660 430868
rect 293132 377692 293188 377702
rect 293244 430388 293300 430398
rect 291564 285172 291620 285182
rect 293132 343140 293188 343150
rect 291452 15922 291508 15932
rect 289772 5954 289828 5964
rect 293132 5908 293188 343084
rect 293244 332578 293300 430332
rect 294924 430164 294980 430174
rect 294812 425458 294868 425468
rect 294812 348598 294868 425402
rect 294924 360298 294980 430108
rect 295260 427588 295316 427598
rect 295036 427476 295092 427486
rect 295036 368758 295092 427420
rect 295260 373798 295316 427532
rect 295260 373732 295316 373742
rect 296492 427252 296548 427262
rect 295036 368692 295092 368702
rect 294924 360232 294980 360242
rect 294812 348532 294868 348542
rect 296492 345178 296548 427196
rect 296604 377578 296660 430802
rect 298284 430500 298340 430510
rect 298172 430138 298228 430148
rect 298060 426898 298116 426908
rect 298060 399700 298116 426842
rect 298060 399634 298116 399644
rect 298172 398020 298228 430082
rect 298172 397954 298228 397964
rect 296604 377512 296660 377522
rect 296492 345112 296548 345122
rect 293244 332512 293300 332522
rect 298172 339108 298228 339118
rect 296492 321636 296548 321646
rect 294812 317604 294868 317614
rect 293244 314218 293300 314228
rect 293244 292292 293300 314162
rect 293244 292226 293300 292236
rect 293132 5842 293188 5852
rect 288092 5058 288148 5068
rect 294812 5124 294868 317548
rect 296492 7588 296548 321580
rect 298172 14308 298228 339052
rect 298284 337438 298340 430444
rect 298396 402778 298452 436156
rect 300748 432964 300804 432974
rect 299964 431038 300020 431048
rect 298620 430276 298676 430286
rect 298396 402712 298452 402722
rect 298508 428518 298564 428528
rect 298508 399588 298564 428462
rect 298620 404578 298676 430220
rect 298620 404512 298676 404522
rect 298732 429604 298788 429614
rect 298508 399522 298564 399532
rect 298732 398098 298788 429548
rect 298956 428484 299012 428494
rect 298956 399476 299012 428428
rect 298956 399410 299012 399420
rect 299852 425098 299908 425108
rect 298732 398032 298788 398042
rect 298284 337372 298340 337382
rect 299852 332398 299908 425042
rect 299852 332332 299908 332342
rect 298172 14242 298228 14252
rect 299852 320292 299908 320302
rect 296492 7522 296548 7532
rect 299852 6020 299908 320236
rect 299964 127558 300020 430982
rect 300748 402388 300804 432908
rect 300860 431060 300916 431070
rect 300860 427438 300916 431004
rect 301084 430948 301140 430958
rect 301084 430678 301140 430892
rect 301084 430622 301812 430678
rect 300860 427372 300916 427382
rect 300972 429940 301028 429950
rect 300748 402322 300804 402332
rect 300860 427140 300916 427150
rect 300860 340138 300916 427084
rect 300972 427078 301028 429884
rect 301084 427922 301700 427978
rect 301084 427812 301140 427922
rect 301084 427746 301140 427756
rect 301532 427438 301588 427448
rect 300972 427022 301140 427078
rect 300972 425278 301028 425288
rect 300972 380436 301028 425222
rect 300972 380370 301028 380380
rect 301084 340318 301140 427022
rect 301532 400596 301588 427382
rect 301644 400708 301700 427922
rect 301756 402724 301812 430622
rect 303212 404398 303268 472562
rect 304448 472350 304768 472384
rect 304448 472294 304518 472350
rect 304574 472294 304642 472350
rect 304698 472294 304768 472350
rect 304448 472226 304768 472294
rect 304448 472170 304518 472226
rect 304574 472170 304642 472226
rect 304698 472170 304768 472226
rect 304448 472102 304768 472170
rect 304448 472046 304518 472102
rect 304574 472046 304642 472102
rect 304698 472046 304768 472102
rect 304448 471978 304768 472046
rect 304448 471922 304518 471978
rect 304574 471922 304642 471978
rect 304698 471922 304768 471978
rect 304448 471888 304768 471922
rect 335168 472350 335488 472384
rect 335168 472294 335238 472350
rect 335294 472294 335362 472350
rect 335418 472294 335488 472350
rect 335168 472226 335488 472294
rect 335168 472170 335238 472226
rect 335294 472170 335362 472226
rect 335418 472170 335488 472226
rect 335168 472102 335488 472170
rect 335168 472046 335238 472102
rect 335294 472046 335362 472102
rect 335418 472046 335488 472102
rect 335168 471978 335488 472046
rect 335168 471922 335238 471978
rect 335294 471922 335362 471978
rect 335418 471922 335488 471978
rect 335168 471888 335488 471922
rect 365888 472350 366208 472384
rect 365888 472294 365958 472350
rect 366014 472294 366082 472350
rect 366138 472294 366208 472350
rect 365888 472226 366208 472294
rect 365888 472170 365958 472226
rect 366014 472170 366082 472226
rect 366138 472170 366208 472226
rect 365888 472102 366208 472170
rect 365888 472046 365958 472102
rect 366014 472046 366082 472102
rect 366138 472046 366208 472102
rect 365888 471978 366208 472046
rect 365888 471922 365958 471978
rect 366014 471922 366082 471978
rect 366138 471922 366208 471978
rect 365888 471888 366208 471922
rect 396608 472350 396928 472384
rect 396608 472294 396678 472350
rect 396734 472294 396802 472350
rect 396858 472294 396928 472350
rect 396608 472226 396928 472294
rect 396608 472170 396678 472226
rect 396734 472170 396802 472226
rect 396858 472170 396928 472226
rect 396608 472102 396928 472170
rect 396608 472046 396678 472102
rect 396734 472046 396802 472102
rect 396858 472046 396928 472102
rect 396608 471978 396928 472046
rect 396608 471922 396678 471978
rect 396734 471922 396802 471978
rect 396858 471922 396928 471978
rect 396608 471888 396928 471922
rect 427328 472350 427648 472384
rect 427328 472294 427398 472350
rect 427454 472294 427522 472350
rect 427578 472294 427648 472350
rect 427328 472226 427648 472294
rect 427328 472170 427398 472226
rect 427454 472170 427522 472226
rect 427578 472170 427648 472226
rect 427328 472102 427648 472170
rect 427328 472046 427398 472102
rect 427454 472046 427522 472102
rect 427578 472046 427648 472102
rect 427328 471978 427648 472046
rect 427328 471922 427398 471978
rect 427454 471922 427522 471978
rect 427578 471922 427648 471978
rect 427328 471888 427648 471922
rect 319808 460350 320128 460384
rect 319808 460294 319878 460350
rect 319934 460294 320002 460350
rect 320058 460294 320128 460350
rect 319808 460226 320128 460294
rect 319808 460170 319878 460226
rect 319934 460170 320002 460226
rect 320058 460170 320128 460226
rect 319808 460102 320128 460170
rect 319808 460046 319878 460102
rect 319934 460046 320002 460102
rect 320058 460046 320128 460102
rect 319808 459978 320128 460046
rect 319808 459922 319878 459978
rect 319934 459922 320002 459978
rect 320058 459922 320128 459978
rect 319808 459888 320128 459922
rect 350528 460350 350848 460384
rect 350528 460294 350598 460350
rect 350654 460294 350722 460350
rect 350778 460294 350848 460350
rect 350528 460226 350848 460294
rect 350528 460170 350598 460226
rect 350654 460170 350722 460226
rect 350778 460170 350848 460226
rect 350528 460102 350848 460170
rect 350528 460046 350598 460102
rect 350654 460046 350722 460102
rect 350778 460046 350848 460102
rect 350528 459978 350848 460046
rect 350528 459922 350598 459978
rect 350654 459922 350722 459978
rect 350778 459922 350848 459978
rect 350528 459888 350848 459922
rect 381248 460350 381568 460384
rect 381248 460294 381318 460350
rect 381374 460294 381442 460350
rect 381498 460294 381568 460350
rect 381248 460226 381568 460294
rect 381248 460170 381318 460226
rect 381374 460170 381442 460226
rect 381498 460170 381568 460226
rect 381248 460102 381568 460170
rect 381248 460046 381318 460102
rect 381374 460046 381442 460102
rect 381498 460046 381568 460102
rect 381248 459978 381568 460046
rect 381248 459922 381318 459978
rect 381374 459922 381442 459978
rect 381498 459922 381568 459978
rect 381248 459888 381568 459922
rect 411968 460350 412288 460384
rect 411968 460294 412038 460350
rect 412094 460294 412162 460350
rect 412218 460294 412288 460350
rect 411968 460226 412288 460294
rect 411968 460170 412038 460226
rect 412094 460170 412162 460226
rect 412218 460170 412288 460226
rect 411968 460102 412288 460170
rect 411968 460046 412038 460102
rect 412094 460046 412162 460102
rect 412218 460046 412288 460102
rect 411968 459978 412288 460046
rect 411968 459922 412038 459978
rect 412094 459922 412162 459978
rect 412218 459922 412288 459978
rect 411968 459888 412288 459922
rect 442688 460350 443008 460384
rect 442688 460294 442758 460350
rect 442814 460294 442882 460350
rect 442938 460294 443008 460350
rect 442688 460226 443008 460294
rect 442688 460170 442758 460226
rect 442814 460170 442882 460226
rect 442938 460170 443008 460226
rect 442688 460102 443008 460170
rect 442688 460046 442758 460102
rect 442814 460046 442882 460102
rect 442938 460046 443008 460102
rect 442688 459978 443008 460046
rect 442688 459922 442758 459978
rect 442814 459922 442882 459978
rect 442938 459922 443008 459978
rect 442688 459888 443008 459922
rect 304448 454350 304768 454384
rect 304448 454294 304518 454350
rect 304574 454294 304642 454350
rect 304698 454294 304768 454350
rect 304448 454226 304768 454294
rect 304448 454170 304518 454226
rect 304574 454170 304642 454226
rect 304698 454170 304768 454226
rect 304448 454102 304768 454170
rect 304448 454046 304518 454102
rect 304574 454046 304642 454102
rect 304698 454046 304768 454102
rect 304448 453978 304768 454046
rect 304448 453922 304518 453978
rect 304574 453922 304642 453978
rect 304698 453922 304768 453978
rect 304448 453888 304768 453922
rect 335168 454350 335488 454384
rect 335168 454294 335238 454350
rect 335294 454294 335362 454350
rect 335418 454294 335488 454350
rect 335168 454226 335488 454294
rect 335168 454170 335238 454226
rect 335294 454170 335362 454226
rect 335418 454170 335488 454226
rect 335168 454102 335488 454170
rect 335168 454046 335238 454102
rect 335294 454046 335362 454102
rect 335418 454046 335488 454102
rect 335168 453978 335488 454046
rect 335168 453922 335238 453978
rect 335294 453922 335362 453978
rect 335418 453922 335488 453978
rect 335168 453888 335488 453922
rect 365888 454350 366208 454384
rect 365888 454294 365958 454350
rect 366014 454294 366082 454350
rect 366138 454294 366208 454350
rect 365888 454226 366208 454294
rect 365888 454170 365958 454226
rect 366014 454170 366082 454226
rect 366138 454170 366208 454226
rect 365888 454102 366208 454170
rect 365888 454046 365958 454102
rect 366014 454046 366082 454102
rect 366138 454046 366208 454102
rect 365888 453978 366208 454046
rect 365888 453922 365958 453978
rect 366014 453922 366082 453978
rect 366138 453922 366208 453978
rect 365888 453888 366208 453922
rect 396608 454350 396928 454384
rect 396608 454294 396678 454350
rect 396734 454294 396802 454350
rect 396858 454294 396928 454350
rect 396608 454226 396928 454294
rect 396608 454170 396678 454226
rect 396734 454170 396802 454226
rect 396858 454170 396928 454226
rect 396608 454102 396928 454170
rect 396608 454046 396678 454102
rect 396734 454046 396802 454102
rect 396858 454046 396928 454102
rect 396608 453978 396928 454046
rect 396608 453922 396678 453978
rect 396734 453922 396802 453978
rect 396858 453922 396928 453978
rect 396608 453888 396928 453922
rect 427328 454350 427648 454384
rect 427328 454294 427398 454350
rect 427454 454294 427522 454350
rect 427578 454294 427648 454350
rect 427328 454226 427648 454294
rect 427328 454170 427398 454226
rect 427454 454170 427522 454226
rect 427578 454170 427648 454226
rect 427328 454102 427648 454170
rect 427328 454046 427398 454102
rect 427454 454046 427522 454102
rect 427578 454046 427648 454102
rect 427328 453978 427648 454046
rect 427328 453922 427398 453978
rect 427454 453922 427522 453978
rect 427578 453922 427648 453978
rect 427328 453888 427648 453922
rect 319808 442350 320128 442384
rect 319808 442294 319878 442350
rect 319934 442294 320002 442350
rect 320058 442294 320128 442350
rect 319808 442226 320128 442294
rect 319808 442170 319878 442226
rect 319934 442170 320002 442226
rect 320058 442170 320128 442226
rect 319808 442102 320128 442170
rect 319808 442046 319878 442102
rect 319934 442046 320002 442102
rect 320058 442046 320128 442102
rect 319808 441978 320128 442046
rect 319808 441922 319878 441978
rect 319934 441922 320002 441978
rect 320058 441922 320128 441978
rect 319808 441888 320128 441922
rect 350528 442350 350848 442384
rect 350528 442294 350598 442350
rect 350654 442294 350722 442350
rect 350778 442294 350848 442350
rect 350528 442226 350848 442294
rect 350528 442170 350598 442226
rect 350654 442170 350722 442226
rect 350778 442170 350848 442226
rect 350528 442102 350848 442170
rect 350528 442046 350598 442102
rect 350654 442046 350722 442102
rect 350778 442046 350848 442102
rect 350528 441978 350848 442046
rect 350528 441922 350598 441978
rect 350654 441922 350722 441978
rect 350778 441922 350848 441978
rect 350528 441888 350848 441922
rect 381248 442350 381568 442384
rect 381248 442294 381318 442350
rect 381374 442294 381442 442350
rect 381498 442294 381568 442350
rect 381248 442226 381568 442294
rect 381248 442170 381318 442226
rect 381374 442170 381442 442226
rect 381498 442170 381568 442226
rect 381248 442102 381568 442170
rect 381248 442046 381318 442102
rect 381374 442046 381442 442102
rect 381498 442046 381568 442102
rect 381248 441978 381568 442046
rect 381248 441922 381318 441978
rect 381374 441922 381442 441978
rect 381498 441922 381568 441978
rect 381248 441888 381568 441922
rect 411968 442350 412288 442384
rect 411968 442294 412038 442350
rect 412094 442294 412162 442350
rect 412218 442294 412288 442350
rect 411968 442226 412288 442294
rect 411968 442170 412038 442226
rect 412094 442170 412162 442226
rect 412218 442170 412288 442226
rect 411968 442102 412288 442170
rect 411968 442046 412038 442102
rect 412094 442046 412162 442102
rect 412218 442046 412288 442102
rect 411968 441978 412288 442046
rect 411968 441922 412038 441978
rect 412094 441922 412162 441978
rect 412218 441922 412288 441978
rect 411968 441888 412288 441922
rect 442688 442350 443008 442384
rect 442688 442294 442758 442350
rect 442814 442294 442882 442350
rect 442938 442294 443008 442350
rect 442688 442226 443008 442294
rect 442688 442170 442758 442226
rect 442814 442170 442882 442226
rect 442938 442170 443008 442226
rect 442688 442102 443008 442170
rect 442688 442046 442758 442102
rect 442814 442046 442882 442102
rect 442938 442046 443008 442102
rect 442688 441978 443008 442046
rect 442688 441922 442758 441978
rect 442814 441922 442882 441978
rect 442938 441922 443008 441978
rect 442688 441888 443008 441922
rect 304448 436350 304768 436384
rect 304448 436294 304518 436350
rect 304574 436294 304642 436350
rect 304698 436294 304768 436350
rect 304448 436226 304768 436294
rect 304448 436170 304518 436226
rect 304574 436170 304642 436226
rect 304698 436170 304768 436226
rect 304448 436102 304768 436170
rect 304448 436046 304518 436102
rect 304574 436046 304642 436102
rect 304698 436046 304768 436102
rect 304448 435978 304768 436046
rect 304448 435922 304518 435978
rect 304574 435922 304642 435978
rect 304698 435922 304768 435978
rect 304448 435888 304768 435922
rect 335168 436350 335488 436384
rect 335168 436294 335238 436350
rect 335294 436294 335362 436350
rect 335418 436294 335488 436350
rect 335168 436226 335488 436294
rect 335168 436170 335238 436226
rect 335294 436170 335362 436226
rect 335418 436170 335488 436226
rect 335168 436102 335488 436170
rect 335168 436046 335238 436102
rect 335294 436046 335362 436102
rect 335418 436046 335488 436102
rect 335168 435978 335488 436046
rect 335168 435922 335238 435978
rect 335294 435922 335362 435978
rect 335418 435922 335488 435978
rect 335168 435888 335488 435922
rect 365888 436350 366208 436384
rect 365888 436294 365958 436350
rect 366014 436294 366082 436350
rect 366138 436294 366208 436350
rect 365888 436226 366208 436294
rect 365888 436170 365958 436226
rect 366014 436170 366082 436226
rect 366138 436170 366208 436226
rect 365888 436102 366208 436170
rect 365888 436046 365958 436102
rect 366014 436046 366082 436102
rect 366138 436046 366208 436102
rect 365888 435978 366208 436046
rect 365888 435922 365958 435978
rect 366014 435922 366082 435978
rect 366138 435922 366208 435978
rect 365888 435888 366208 435922
rect 396608 436350 396928 436384
rect 396608 436294 396678 436350
rect 396734 436294 396802 436350
rect 396858 436294 396928 436350
rect 396608 436226 396928 436294
rect 396608 436170 396678 436226
rect 396734 436170 396802 436226
rect 396858 436170 396928 436226
rect 396608 436102 396928 436170
rect 396608 436046 396678 436102
rect 396734 436046 396802 436102
rect 396858 436046 396928 436102
rect 396608 435978 396928 436046
rect 396608 435922 396678 435978
rect 396734 435922 396802 435978
rect 396858 435922 396928 435978
rect 396608 435888 396928 435922
rect 427328 436350 427648 436384
rect 427328 436294 427398 436350
rect 427454 436294 427522 436350
rect 427578 436294 427648 436350
rect 427328 436226 427648 436294
rect 427328 436170 427398 436226
rect 427454 436170 427522 436226
rect 427578 436170 427648 436226
rect 427328 436102 427648 436170
rect 427328 436046 427398 436102
rect 427454 436046 427522 436102
rect 427578 436046 427648 436102
rect 427328 435978 427648 436046
rect 427328 435922 427398 435978
rect 427454 435922 427522 435978
rect 427578 435922 427648 435978
rect 427328 435888 427648 435922
rect 452732 433378 452788 551222
rect 452732 433312 452788 433322
rect 457772 548218 457828 548228
rect 457772 432628 457828 548162
rect 457772 432562 457828 432572
rect 319808 424350 320128 424384
rect 319808 424294 319878 424350
rect 319934 424294 320002 424350
rect 320058 424294 320128 424350
rect 319808 424226 320128 424294
rect 319808 424170 319878 424226
rect 319934 424170 320002 424226
rect 320058 424170 320128 424226
rect 319808 424102 320128 424170
rect 319808 424046 319878 424102
rect 319934 424046 320002 424102
rect 320058 424046 320128 424102
rect 319808 423978 320128 424046
rect 319808 423922 319878 423978
rect 319934 423922 320002 423978
rect 320058 423922 320128 423978
rect 319808 423888 320128 423922
rect 350528 424350 350848 424384
rect 350528 424294 350598 424350
rect 350654 424294 350722 424350
rect 350778 424294 350848 424350
rect 350528 424226 350848 424294
rect 350528 424170 350598 424226
rect 350654 424170 350722 424226
rect 350778 424170 350848 424226
rect 350528 424102 350848 424170
rect 350528 424046 350598 424102
rect 350654 424046 350722 424102
rect 350778 424046 350848 424102
rect 350528 423978 350848 424046
rect 350528 423922 350598 423978
rect 350654 423922 350722 423978
rect 350778 423922 350848 423978
rect 350528 423888 350848 423922
rect 381248 424350 381568 424384
rect 381248 424294 381318 424350
rect 381374 424294 381442 424350
rect 381498 424294 381568 424350
rect 381248 424226 381568 424294
rect 381248 424170 381318 424226
rect 381374 424170 381442 424226
rect 381498 424170 381568 424226
rect 381248 424102 381568 424170
rect 381248 424046 381318 424102
rect 381374 424046 381442 424102
rect 381498 424046 381568 424102
rect 381248 423978 381568 424046
rect 381248 423922 381318 423978
rect 381374 423922 381442 423978
rect 381498 423922 381568 423978
rect 381248 423888 381568 423922
rect 411968 424350 412288 424384
rect 411968 424294 412038 424350
rect 412094 424294 412162 424350
rect 412218 424294 412288 424350
rect 411968 424226 412288 424294
rect 411968 424170 412038 424226
rect 412094 424170 412162 424226
rect 412218 424170 412288 424226
rect 411968 424102 412288 424170
rect 411968 424046 412038 424102
rect 412094 424046 412162 424102
rect 412218 424046 412288 424102
rect 411968 423978 412288 424046
rect 411968 423922 412038 423978
rect 412094 423922 412162 423978
rect 412218 423922 412288 423978
rect 411968 423888 412288 423922
rect 442688 424350 443008 424384
rect 442688 424294 442758 424350
rect 442814 424294 442882 424350
rect 442938 424294 443008 424350
rect 442688 424226 443008 424294
rect 442688 424170 442758 424226
rect 442814 424170 442882 424226
rect 442938 424170 443008 424226
rect 442688 424102 443008 424170
rect 442688 424046 442758 424102
rect 442814 424046 442882 424102
rect 442938 424046 443008 424102
rect 442688 423978 443008 424046
rect 442688 423922 442758 423978
rect 442814 423922 442882 423978
rect 442938 423922 443008 423978
rect 442688 423888 443008 423922
rect 304448 418350 304768 418384
rect 304448 418294 304518 418350
rect 304574 418294 304642 418350
rect 304698 418294 304768 418350
rect 304448 418226 304768 418294
rect 304448 418170 304518 418226
rect 304574 418170 304642 418226
rect 304698 418170 304768 418226
rect 304448 418102 304768 418170
rect 304448 418046 304518 418102
rect 304574 418046 304642 418102
rect 304698 418046 304768 418102
rect 304448 417978 304768 418046
rect 304448 417922 304518 417978
rect 304574 417922 304642 417978
rect 304698 417922 304768 417978
rect 304448 417888 304768 417922
rect 335168 418350 335488 418384
rect 335168 418294 335238 418350
rect 335294 418294 335362 418350
rect 335418 418294 335488 418350
rect 335168 418226 335488 418294
rect 335168 418170 335238 418226
rect 335294 418170 335362 418226
rect 335418 418170 335488 418226
rect 335168 418102 335488 418170
rect 335168 418046 335238 418102
rect 335294 418046 335362 418102
rect 335418 418046 335488 418102
rect 335168 417978 335488 418046
rect 335168 417922 335238 417978
rect 335294 417922 335362 417978
rect 335418 417922 335488 417978
rect 335168 417888 335488 417922
rect 365888 418350 366208 418384
rect 365888 418294 365958 418350
rect 366014 418294 366082 418350
rect 366138 418294 366208 418350
rect 365888 418226 366208 418294
rect 365888 418170 365958 418226
rect 366014 418170 366082 418226
rect 366138 418170 366208 418226
rect 365888 418102 366208 418170
rect 365888 418046 365958 418102
rect 366014 418046 366082 418102
rect 366138 418046 366208 418102
rect 365888 417978 366208 418046
rect 365888 417922 365958 417978
rect 366014 417922 366082 417978
rect 366138 417922 366208 417978
rect 365888 417888 366208 417922
rect 396608 418350 396928 418384
rect 396608 418294 396678 418350
rect 396734 418294 396802 418350
rect 396858 418294 396928 418350
rect 396608 418226 396928 418294
rect 396608 418170 396678 418226
rect 396734 418170 396802 418226
rect 396858 418170 396928 418226
rect 396608 418102 396928 418170
rect 396608 418046 396678 418102
rect 396734 418046 396802 418102
rect 396858 418046 396928 418102
rect 396608 417978 396928 418046
rect 396608 417922 396678 417978
rect 396734 417922 396802 417978
rect 396858 417922 396928 417978
rect 396608 417888 396928 417922
rect 427328 418350 427648 418384
rect 427328 418294 427398 418350
rect 427454 418294 427522 418350
rect 427578 418294 427648 418350
rect 427328 418226 427648 418294
rect 427328 418170 427398 418226
rect 427454 418170 427522 418226
rect 427578 418170 427648 418226
rect 427328 418102 427648 418170
rect 427328 418046 427398 418102
rect 427454 418046 427522 418102
rect 427578 418046 427648 418102
rect 427328 417978 427648 418046
rect 427328 417922 427398 417978
rect 427454 417922 427522 417978
rect 427578 417922 427648 417978
rect 427328 417888 427648 417922
rect 451052 411908 451108 411918
rect 449372 410340 449428 410350
rect 319808 406350 320128 406384
rect 319808 406294 319878 406350
rect 319934 406294 320002 406350
rect 320058 406294 320128 406350
rect 319808 406226 320128 406294
rect 319808 406170 319878 406226
rect 319934 406170 320002 406226
rect 320058 406170 320128 406226
rect 319808 406102 320128 406170
rect 319808 406046 319878 406102
rect 319934 406046 320002 406102
rect 320058 406046 320128 406102
rect 319808 405978 320128 406046
rect 319808 405922 319878 405978
rect 319934 405922 320002 405978
rect 320058 405922 320128 405978
rect 319808 405888 320128 405922
rect 350528 406350 350848 406384
rect 350528 406294 350598 406350
rect 350654 406294 350722 406350
rect 350778 406294 350848 406350
rect 350528 406226 350848 406294
rect 350528 406170 350598 406226
rect 350654 406170 350722 406226
rect 350778 406170 350848 406226
rect 350528 406102 350848 406170
rect 350528 406046 350598 406102
rect 350654 406046 350722 406102
rect 350778 406046 350848 406102
rect 350528 405978 350848 406046
rect 350528 405922 350598 405978
rect 350654 405922 350722 405978
rect 350778 405922 350848 405978
rect 350528 405888 350848 405922
rect 381248 406350 381568 406384
rect 381248 406294 381318 406350
rect 381374 406294 381442 406350
rect 381498 406294 381568 406350
rect 381248 406226 381568 406294
rect 381248 406170 381318 406226
rect 381374 406170 381442 406226
rect 381498 406170 381568 406226
rect 381248 406102 381568 406170
rect 381248 406046 381318 406102
rect 381374 406046 381442 406102
rect 381498 406046 381568 406102
rect 381248 405978 381568 406046
rect 381248 405922 381318 405978
rect 381374 405922 381442 405978
rect 381498 405922 381568 405978
rect 381248 405888 381568 405922
rect 411968 406350 412288 406384
rect 411968 406294 412038 406350
rect 412094 406294 412162 406350
rect 412218 406294 412288 406350
rect 411968 406226 412288 406294
rect 411968 406170 412038 406226
rect 412094 406170 412162 406226
rect 412218 406170 412288 406226
rect 411968 406102 412288 406170
rect 411968 406046 412038 406102
rect 412094 406046 412162 406102
rect 412218 406046 412288 406102
rect 411968 405978 412288 406046
rect 411968 405922 412038 405978
rect 412094 405922 412162 405978
rect 412218 405922 412288 405978
rect 411968 405888 412288 405922
rect 442688 406350 443008 406384
rect 442688 406294 442758 406350
rect 442814 406294 442882 406350
rect 442938 406294 443008 406350
rect 442688 406226 443008 406294
rect 442688 406170 442758 406226
rect 442814 406170 442882 406226
rect 442938 406170 443008 406226
rect 442688 406102 443008 406170
rect 442688 406046 442758 406102
rect 442814 406046 442882 406102
rect 442938 406046 443008 406102
rect 442688 405978 443008 406046
rect 442688 405922 442758 405978
rect 442814 405922 442882 405978
rect 442938 405922 443008 405978
rect 442688 405888 443008 405922
rect 303212 404332 303268 404342
rect 301756 402658 301812 402668
rect 301644 400642 301700 400652
rect 301532 400530 301588 400540
rect 312618 400350 313238 402722
rect 312618 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 313238 400350
rect 312618 400226 313238 400294
rect 312618 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 313238 400226
rect 312618 400102 313238 400170
rect 312618 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 313238 400102
rect 312618 399978 313238 400046
rect 312618 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 313238 399978
rect 312618 382350 313238 399922
rect 312618 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 313238 382350
rect 312618 382226 313238 382294
rect 312618 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 313238 382226
rect 312618 382102 313238 382170
rect 312618 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 313238 382102
rect 312618 381978 313238 382046
rect 312618 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 313238 381978
rect 301908 370350 302384 370384
rect 301908 370294 301932 370350
rect 301988 370294 302056 370350
rect 302112 370294 302180 370350
rect 302236 370294 302304 370350
rect 302360 370294 302384 370350
rect 301908 370226 302384 370294
rect 301908 370170 301932 370226
rect 301988 370170 302056 370226
rect 302112 370170 302180 370226
rect 302236 370170 302304 370226
rect 302360 370170 302384 370226
rect 301908 370102 302384 370170
rect 301908 370046 301932 370102
rect 301988 370046 302056 370102
rect 302112 370046 302180 370102
rect 302236 370046 302304 370102
rect 302360 370046 302384 370102
rect 301908 369978 302384 370046
rect 301908 369922 301932 369978
rect 301988 369922 302056 369978
rect 302112 369922 302180 369978
rect 302236 369922 302304 369978
rect 302360 369922 302384 369978
rect 301908 369888 302384 369922
rect 302708 364350 303184 364384
rect 302708 364294 302732 364350
rect 302788 364294 302856 364350
rect 302912 364294 302980 364350
rect 303036 364294 303104 364350
rect 303160 364294 303184 364350
rect 302708 364226 303184 364294
rect 302708 364170 302732 364226
rect 302788 364170 302856 364226
rect 302912 364170 302980 364226
rect 303036 364170 303104 364226
rect 303160 364170 303184 364226
rect 302708 364102 303184 364170
rect 302708 364046 302732 364102
rect 302788 364046 302856 364102
rect 302912 364046 302980 364102
rect 303036 364046 303104 364102
rect 303160 364046 303184 364102
rect 302708 363978 303184 364046
rect 302708 363922 302732 363978
rect 302788 363922 302856 363978
rect 302912 363922 302980 363978
rect 303036 363922 303104 363978
rect 303160 363922 303184 363978
rect 302708 363888 303184 363922
rect 312618 364350 313238 381922
rect 312618 364294 312714 364350
rect 312770 364294 312838 364350
rect 312894 364294 312962 364350
rect 313018 364294 313086 364350
rect 313142 364294 313238 364350
rect 312618 364226 313238 364294
rect 312618 364170 312714 364226
rect 312770 364170 312838 364226
rect 312894 364170 312962 364226
rect 313018 364170 313086 364226
rect 313142 364170 313238 364226
rect 312618 364102 313238 364170
rect 312618 364046 312714 364102
rect 312770 364046 312838 364102
rect 312894 364046 312962 364102
rect 313018 364046 313086 364102
rect 313142 364046 313238 364102
rect 312618 363978 313238 364046
rect 312618 363922 312714 363978
rect 312770 363922 312838 363978
rect 312894 363922 312962 363978
rect 313018 363922 313086 363978
rect 313142 363922 313238 363978
rect 301908 352350 302384 352384
rect 301908 352294 301932 352350
rect 301988 352294 302056 352350
rect 302112 352294 302180 352350
rect 302236 352294 302304 352350
rect 302360 352294 302384 352350
rect 301908 352226 302384 352294
rect 301908 352170 301932 352226
rect 301988 352170 302056 352226
rect 302112 352170 302180 352226
rect 302236 352170 302304 352226
rect 302360 352170 302384 352226
rect 301908 352102 302384 352170
rect 301908 352046 301932 352102
rect 301988 352046 302056 352102
rect 302112 352046 302180 352102
rect 302236 352046 302304 352102
rect 302360 352046 302384 352102
rect 301908 351978 302384 352046
rect 301908 351922 301932 351978
rect 301988 351922 302056 351978
rect 302112 351922 302180 351978
rect 302236 351922 302304 351978
rect 302360 351922 302384 351978
rect 301908 351888 302384 351922
rect 302708 346350 303184 346384
rect 302708 346294 302732 346350
rect 302788 346294 302856 346350
rect 302912 346294 302980 346350
rect 303036 346294 303104 346350
rect 303160 346294 303184 346350
rect 302708 346226 303184 346294
rect 302708 346170 302732 346226
rect 302788 346170 302856 346226
rect 302912 346170 302980 346226
rect 303036 346170 303104 346226
rect 303160 346170 303184 346226
rect 302708 346102 303184 346170
rect 302708 346046 302732 346102
rect 302788 346046 302856 346102
rect 302912 346046 302980 346102
rect 303036 346046 303104 346102
rect 303160 346046 303184 346102
rect 302708 345978 303184 346046
rect 302708 345922 302732 345978
rect 302788 345922 302856 345978
rect 302912 345922 302980 345978
rect 303036 345922 303104 345978
rect 303160 345922 303184 345978
rect 302708 345888 303184 345922
rect 312618 346350 313238 363922
rect 312618 346294 312714 346350
rect 312770 346294 312838 346350
rect 312894 346294 312962 346350
rect 313018 346294 313086 346350
rect 313142 346294 313238 346350
rect 312618 346226 313238 346294
rect 312618 346170 312714 346226
rect 312770 346170 312838 346226
rect 312894 346170 312962 346226
rect 313018 346170 313086 346226
rect 313142 346170 313238 346226
rect 312618 346102 313238 346170
rect 312618 346046 312714 346102
rect 312770 346046 312838 346102
rect 312894 346046 312962 346102
rect 313018 346046 313086 346102
rect 313142 346046 313238 346102
rect 312618 345978 313238 346046
rect 312618 345922 312714 345978
rect 312770 345922 312838 345978
rect 312894 345922 312962 345978
rect 313018 345922 313086 345978
rect 313142 345922 313238 345978
rect 301084 340252 301140 340262
rect 300860 340072 300916 340082
rect 301908 334350 302384 334384
rect 301908 334294 301932 334350
rect 301988 334294 302056 334350
rect 302112 334294 302180 334350
rect 302236 334294 302304 334350
rect 302360 334294 302384 334350
rect 301908 334226 302384 334294
rect 301908 334170 301932 334226
rect 301988 334170 302056 334226
rect 302112 334170 302180 334226
rect 302236 334170 302304 334226
rect 302360 334170 302384 334226
rect 301908 334102 302384 334170
rect 301908 334046 301932 334102
rect 301988 334046 302056 334102
rect 302112 334046 302180 334102
rect 302236 334046 302304 334102
rect 302360 334046 302384 334102
rect 301908 333978 302384 334046
rect 301908 333922 301932 333978
rect 301988 333922 302056 333978
rect 302112 333922 302180 333978
rect 302236 333922 302304 333978
rect 302360 333922 302384 333978
rect 301908 333888 302384 333922
rect 302708 328350 303184 328384
rect 302708 328294 302732 328350
rect 302788 328294 302856 328350
rect 302912 328294 302980 328350
rect 303036 328294 303104 328350
rect 303160 328294 303184 328350
rect 302708 328226 303184 328294
rect 302708 328170 302732 328226
rect 302788 328170 302856 328226
rect 302912 328170 302980 328226
rect 303036 328170 303104 328226
rect 303160 328170 303184 328226
rect 302708 328102 303184 328170
rect 302708 328046 302732 328102
rect 302788 328046 302856 328102
rect 302912 328046 302980 328102
rect 303036 328046 303104 328102
rect 303160 328046 303184 328102
rect 302708 327978 303184 328046
rect 302708 327922 302732 327978
rect 302788 327922 302856 327978
rect 302912 327922 302980 327978
rect 303036 327922 303104 327978
rect 303160 327922 303184 327978
rect 302708 327888 303184 327922
rect 312618 328350 313238 345922
rect 312618 328294 312714 328350
rect 312770 328294 312838 328350
rect 312894 328294 312962 328350
rect 313018 328294 313086 328350
rect 313142 328294 313238 328350
rect 312618 328226 313238 328294
rect 312618 328170 312714 328226
rect 312770 328170 312838 328226
rect 312894 328170 312962 328226
rect 313018 328170 313086 328226
rect 313142 328170 313238 328226
rect 312618 328102 313238 328170
rect 312618 328046 312714 328102
rect 312770 328046 312838 328102
rect 312894 328046 312962 328102
rect 313018 328046 313086 328102
rect 313142 328046 313238 328102
rect 312618 327978 313238 328046
rect 312618 327922 312714 327978
rect 312770 327922 312838 327978
rect 312894 327922 312962 327978
rect 313018 327922 313086 327978
rect 313142 327922 313238 327978
rect 301908 316350 302384 316384
rect 301908 316294 301932 316350
rect 301988 316294 302056 316350
rect 302112 316294 302180 316350
rect 302236 316294 302304 316350
rect 302360 316294 302384 316350
rect 301908 316226 302384 316294
rect 301908 316170 301932 316226
rect 301988 316170 302056 316226
rect 302112 316170 302180 316226
rect 302236 316170 302304 316226
rect 302360 316170 302384 316226
rect 301908 316102 302384 316170
rect 301908 316046 301932 316102
rect 301988 316046 302056 316102
rect 302112 316046 302180 316102
rect 302236 316046 302304 316102
rect 302360 316046 302384 316102
rect 301908 315978 302384 316046
rect 301908 315922 301932 315978
rect 301988 315922 302056 315978
rect 302112 315922 302180 315978
rect 302236 315922 302304 315978
rect 302360 315922 302384 315978
rect 301908 315888 302384 315922
rect 302708 310350 303184 310384
rect 302708 310294 302732 310350
rect 302788 310294 302856 310350
rect 302912 310294 302980 310350
rect 303036 310294 303104 310350
rect 303160 310294 303184 310350
rect 302708 310226 303184 310294
rect 302708 310170 302732 310226
rect 302788 310170 302856 310226
rect 302912 310170 302980 310226
rect 303036 310170 303104 310226
rect 303160 310170 303184 310226
rect 302708 310102 303184 310170
rect 302708 310046 302732 310102
rect 302788 310046 302856 310102
rect 302912 310046 302980 310102
rect 303036 310046 303104 310102
rect 303160 310046 303184 310102
rect 302708 309978 303184 310046
rect 302708 309922 302732 309978
rect 302788 309922 302856 309978
rect 302912 309922 302980 309978
rect 303036 309922 303104 309978
rect 303160 309922 303184 309978
rect 302708 309888 303184 309922
rect 312618 310350 313238 327922
rect 312618 310294 312714 310350
rect 312770 310294 312838 310350
rect 312894 310294 312962 310350
rect 313018 310294 313086 310350
rect 313142 310294 313238 310350
rect 312618 310226 313238 310294
rect 312618 310170 312714 310226
rect 312770 310170 312838 310226
rect 312894 310170 312962 310226
rect 313018 310170 313086 310226
rect 313142 310170 313238 310226
rect 312618 310102 313238 310170
rect 312618 310046 312714 310102
rect 312770 310046 312838 310102
rect 312894 310046 312962 310102
rect 313018 310046 313086 310102
rect 313142 310046 313238 310102
rect 312618 309978 313238 310046
rect 312618 309922 312714 309978
rect 312770 309922 312838 309978
rect 312894 309922 312962 309978
rect 313018 309922 313086 309978
rect 313142 309922 313238 309978
rect 301908 298350 302384 298384
rect 301908 298294 301932 298350
rect 301988 298294 302056 298350
rect 302112 298294 302180 298350
rect 302236 298294 302304 298350
rect 302360 298294 302384 298350
rect 301908 298226 302384 298294
rect 301908 298170 301932 298226
rect 301988 298170 302056 298226
rect 302112 298170 302180 298226
rect 302236 298170 302304 298226
rect 302360 298170 302384 298226
rect 301908 298102 302384 298170
rect 301908 298046 301932 298102
rect 301988 298046 302056 298102
rect 302112 298046 302180 298102
rect 302236 298046 302304 298102
rect 302360 298046 302384 298102
rect 301908 297978 302384 298046
rect 301908 297922 301932 297978
rect 301988 297922 302056 297978
rect 302112 297922 302180 297978
rect 302236 297922 302304 297978
rect 302360 297922 302384 297978
rect 301908 297888 302384 297922
rect 302708 292350 303184 292384
rect 302708 292294 302732 292350
rect 302788 292294 302856 292350
rect 302912 292294 302980 292350
rect 303036 292294 303104 292350
rect 303160 292294 303184 292350
rect 302708 292226 303184 292294
rect 302708 292170 302732 292226
rect 302788 292170 302856 292226
rect 302912 292170 302980 292226
rect 303036 292170 303104 292226
rect 303160 292170 303184 292226
rect 302708 292102 303184 292170
rect 302708 292046 302732 292102
rect 302788 292046 302856 292102
rect 302912 292046 302980 292102
rect 303036 292046 303104 292102
rect 303160 292046 303184 292102
rect 302708 291978 303184 292046
rect 302708 291922 302732 291978
rect 302788 291922 302856 291978
rect 302912 291922 302980 291978
rect 303036 291922 303104 291978
rect 303160 291922 303184 291978
rect 302708 291888 303184 291922
rect 312618 292350 313238 309922
rect 312618 292294 312714 292350
rect 312770 292294 312838 292350
rect 312894 292294 312962 292350
rect 313018 292294 313086 292350
rect 313142 292294 313238 292350
rect 312618 292226 313238 292294
rect 312618 292170 312714 292226
rect 312770 292170 312838 292226
rect 312894 292170 312962 292226
rect 313018 292170 313086 292226
rect 313142 292170 313238 292226
rect 312618 292102 313238 292170
rect 312618 292046 312714 292102
rect 312770 292046 312838 292102
rect 312894 292046 312962 292102
rect 313018 292046 313086 292102
rect 313142 292046 313238 292102
rect 312618 291978 313238 292046
rect 312618 291922 312714 291978
rect 312770 291922 312838 291978
rect 312894 291922 312962 291978
rect 313018 291922 313086 291978
rect 313142 291922 313238 291978
rect 304892 279972 304948 279982
rect 304780 142772 304836 142782
rect 304780 142138 304836 142716
rect 304780 142072 304836 142082
rect 303996 140878 304052 140888
rect 303996 140644 304052 140822
rect 303996 140578 304052 140588
rect 299964 127492 300020 127502
rect 299852 5954 299908 5964
rect 294812 5058 294868 5068
rect 304892 4228 304948 279916
rect 304892 4162 304948 4172
rect 312618 274350 313238 291922
rect 312618 274294 312714 274350
rect 312770 274294 312838 274350
rect 312894 274294 312962 274350
rect 313018 274294 313086 274350
rect 313142 274294 313238 274350
rect 312618 274226 313238 274294
rect 312618 274170 312714 274226
rect 312770 274170 312838 274226
rect 312894 274170 312962 274226
rect 313018 274170 313086 274226
rect 313142 274170 313238 274226
rect 312618 274102 313238 274170
rect 312618 274046 312714 274102
rect 312770 274046 312838 274102
rect 312894 274046 312962 274102
rect 313018 274046 313086 274102
rect 313142 274046 313238 274102
rect 312618 273978 313238 274046
rect 312618 273922 312714 273978
rect 312770 273922 312838 273978
rect 312894 273922 312962 273978
rect 313018 273922 313086 273978
rect 313142 273922 313238 273978
rect 312618 256350 313238 273922
rect 312618 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 313238 256350
rect 312618 256226 313238 256294
rect 312618 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 313238 256226
rect 312618 256102 313238 256170
rect 312618 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 313238 256102
rect 312618 255978 313238 256046
rect 312618 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 313238 255978
rect 312618 238350 313238 255922
rect 312618 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 313238 238350
rect 312618 238226 313238 238294
rect 312618 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 313238 238226
rect 312618 238102 313238 238170
rect 312618 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 313238 238102
rect 312618 237978 313238 238046
rect 312618 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 313238 237978
rect 312618 220350 313238 237922
rect 312618 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 313238 220350
rect 312618 220226 313238 220294
rect 312618 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 313238 220226
rect 312618 220102 313238 220170
rect 312618 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 313238 220102
rect 312618 219978 313238 220046
rect 312618 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 313238 219978
rect 312618 202350 313238 219922
rect 312618 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 313238 202350
rect 312618 202226 313238 202294
rect 312618 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 313238 202226
rect 312618 202102 313238 202170
rect 312618 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 313238 202102
rect 312618 201978 313238 202046
rect 312618 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 313238 201978
rect 312618 184350 313238 201922
rect 312618 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 313238 184350
rect 312618 184226 313238 184294
rect 312618 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 313238 184226
rect 312618 184102 313238 184170
rect 312618 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 313238 184102
rect 312618 183978 313238 184046
rect 312618 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 313238 183978
rect 312618 166350 313238 183922
rect 312618 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 313238 166350
rect 312618 166226 313238 166294
rect 312618 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 313238 166226
rect 312618 166102 313238 166170
rect 312618 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 313238 166102
rect 312618 165978 313238 166046
rect 312618 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 313238 165978
rect 312618 148350 313238 165922
rect 312618 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 313238 148350
rect 312618 148226 313238 148294
rect 312618 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 313238 148226
rect 312618 148102 313238 148170
rect 312618 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 313238 148102
rect 312618 147978 313238 148046
rect 312618 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 313238 147978
rect 312618 130350 313238 147922
rect 316338 388350 316958 402722
rect 316338 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 316958 388350
rect 316338 388226 316958 388294
rect 316338 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 316958 388226
rect 316338 388102 316958 388170
rect 316338 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 316958 388102
rect 316338 387978 316958 388046
rect 316338 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 316958 387978
rect 316338 370350 316958 387922
rect 316338 370294 316434 370350
rect 316490 370294 316558 370350
rect 316614 370294 316682 370350
rect 316738 370294 316806 370350
rect 316862 370294 316958 370350
rect 316338 370226 316958 370294
rect 316338 370170 316434 370226
rect 316490 370170 316558 370226
rect 316614 370170 316682 370226
rect 316738 370170 316806 370226
rect 316862 370170 316958 370226
rect 316338 370102 316958 370170
rect 316338 370046 316434 370102
rect 316490 370046 316558 370102
rect 316614 370046 316682 370102
rect 316738 370046 316806 370102
rect 316862 370046 316958 370102
rect 316338 369978 316958 370046
rect 316338 369922 316434 369978
rect 316490 369922 316558 369978
rect 316614 369922 316682 369978
rect 316738 369922 316806 369978
rect 316862 369922 316958 369978
rect 316338 352350 316958 369922
rect 316338 352294 316434 352350
rect 316490 352294 316558 352350
rect 316614 352294 316682 352350
rect 316738 352294 316806 352350
rect 316862 352294 316958 352350
rect 316338 352226 316958 352294
rect 316338 352170 316434 352226
rect 316490 352170 316558 352226
rect 316614 352170 316682 352226
rect 316738 352170 316806 352226
rect 316862 352170 316958 352226
rect 316338 352102 316958 352170
rect 316338 352046 316434 352102
rect 316490 352046 316558 352102
rect 316614 352046 316682 352102
rect 316738 352046 316806 352102
rect 316862 352046 316958 352102
rect 316338 351978 316958 352046
rect 316338 351922 316434 351978
rect 316490 351922 316558 351978
rect 316614 351922 316682 351978
rect 316738 351922 316806 351978
rect 316862 351922 316958 351978
rect 316338 334350 316958 351922
rect 316338 334294 316434 334350
rect 316490 334294 316558 334350
rect 316614 334294 316682 334350
rect 316738 334294 316806 334350
rect 316862 334294 316958 334350
rect 316338 334226 316958 334294
rect 316338 334170 316434 334226
rect 316490 334170 316558 334226
rect 316614 334170 316682 334226
rect 316738 334170 316806 334226
rect 316862 334170 316958 334226
rect 316338 334102 316958 334170
rect 316338 334046 316434 334102
rect 316490 334046 316558 334102
rect 316614 334046 316682 334102
rect 316738 334046 316806 334102
rect 316862 334046 316958 334102
rect 316338 333978 316958 334046
rect 316338 333922 316434 333978
rect 316490 333922 316558 333978
rect 316614 333922 316682 333978
rect 316738 333922 316806 333978
rect 316862 333922 316958 333978
rect 316338 316350 316958 333922
rect 316338 316294 316434 316350
rect 316490 316294 316558 316350
rect 316614 316294 316682 316350
rect 316738 316294 316806 316350
rect 316862 316294 316958 316350
rect 316338 316226 316958 316294
rect 316338 316170 316434 316226
rect 316490 316170 316558 316226
rect 316614 316170 316682 316226
rect 316738 316170 316806 316226
rect 316862 316170 316958 316226
rect 316338 316102 316958 316170
rect 316338 316046 316434 316102
rect 316490 316046 316558 316102
rect 316614 316046 316682 316102
rect 316738 316046 316806 316102
rect 316862 316046 316958 316102
rect 316338 315978 316958 316046
rect 316338 315922 316434 315978
rect 316490 315922 316558 315978
rect 316614 315922 316682 315978
rect 316738 315922 316806 315978
rect 316862 315922 316958 315978
rect 316338 298350 316958 315922
rect 316338 298294 316434 298350
rect 316490 298294 316558 298350
rect 316614 298294 316682 298350
rect 316738 298294 316806 298350
rect 316862 298294 316958 298350
rect 316338 298226 316958 298294
rect 316338 298170 316434 298226
rect 316490 298170 316558 298226
rect 316614 298170 316682 298226
rect 316738 298170 316806 298226
rect 316862 298170 316958 298226
rect 316338 298102 316958 298170
rect 316338 298046 316434 298102
rect 316490 298046 316558 298102
rect 316614 298046 316682 298102
rect 316738 298046 316806 298102
rect 316862 298046 316958 298102
rect 316338 297978 316958 298046
rect 316338 297922 316434 297978
rect 316490 297922 316558 297978
rect 316614 297922 316682 297978
rect 316738 297922 316806 297978
rect 316862 297922 316958 297978
rect 316338 280350 316958 297922
rect 316338 280294 316434 280350
rect 316490 280294 316558 280350
rect 316614 280294 316682 280350
rect 316738 280294 316806 280350
rect 316862 280294 316958 280350
rect 316338 280226 316958 280294
rect 316338 280170 316434 280226
rect 316490 280170 316558 280226
rect 316614 280170 316682 280226
rect 316738 280170 316806 280226
rect 316862 280170 316958 280226
rect 316338 280102 316958 280170
rect 316338 280046 316434 280102
rect 316490 280046 316558 280102
rect 316614 280046 316682 280102
rect 316738 280046 316806 280102
rect 316862 280046 316958 280102
rect 316338 279978 316958 280046
rect 316338 279922 316434 279978
rect 316490 279922 316558 279978
rect 316614 279922 316682 279978
rect 316738 279922 316806 279978
rect 316862 279922 316958 279978
rect 316338 262350 316958 279922
rect 316338 262294 316434 262350
rect 316490 262294 316558 262350
rect 316614 262294 316682 262350
rect 316738 262294 316806 262350
rect 316862 262294 316958 262350
rect 316338 262226 316958 262294
rect 316338 262170 316434 262226
rect 316490 262170 316558 262226
rect 316614 262170 316682 262226
rect 316738 262170 316806 262226
rect 316862 262170 316958 262226
rect 316338 262102 316958 262170
rect 316338 262046 316434 262102
rect 316490 262046 316558 262102
rect 316614 262046 316682 262102
rect 316738 262046 316806 262102
rect 316862 262046 316958 262102
rect 316338 261978 316958 262046
rect 316338 261922 316434 261978
rect 316490 261922 316558 261978
rect 316614 261922 316682 261978
rect 316738 261922 316806 261978
rect 316862 261922 316958 261978
rect 316338 244350 316958 261922
rect 316338 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 316958 244350
rect 316338 244226 316958 244294
rect 316338 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 316958 244226
rect 316338 244102 316958 244170
rect 316338 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 316958 244102
rect 316338 243978 316958 244046
rect 316338 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 316958 243978
rect 316338 226350 316958 243922
rect 316338 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 316958 226350
rect 316338 226226 316958 226294
rect 316338 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 316958 226226
rect 316338 226102 316958 226170
rect 316338 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 316958 226102
rect 316338 225978 316958 226046
rect 316338 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 316958 225978
rect 316338 208350 316958 225922
rect 316338 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 316958 208350
rect 316338 208226 316958 208294
rect 316338 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 316958 208226
rect 316338 208102 316958 208170
rect 316338 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 316958 208102
rect 316338 207978 316958 208046
rect 316338 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 316958 207978
rect 316338 190350 316958 207922
rect 316338 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 316958 190350
rect 316338 190226 316958 190294
rect 316338 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 316958 190226
rect 316338 190102 316958 190170
rect 316338 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 316958 190102
rect 316338 189978 316958 190046
rect 316338 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 316958 189978
rect 316338 172350 316958 189922
rect 316338 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 316958 172350
rect 316338 172226 316958 172294
rect 316338 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 316958 172226
rect 316338 172102 316958 172170
rect 316338 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 316958 172102
rect 316338 171978 316958 172046
rect 316338 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 316958 171978
rect 316338 154350 316958 171922
rect 343338 400350 343958 402722
rect 343338 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 343958 400350
rect 343338 400226 343958 400294
rect 343338 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 343958 400226
rect 343338 400102 343958 400170
rect 343338 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 343958 400102
rect 343338 399978 343958 400046
rect 343338 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 343958 399978
rect 343338 382350 343958 399922
rect 343338 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 343958 382350
rect 343338 382226 343958 382294
rect 343338 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 343958 382226
rect 343338 382102 343958 382170
rect 343338 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 343958 382102
rect 343338 381978 343958 382046
rect 343338 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 343958 381978
rect 343338 364350 343958 381922
rect 343338 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 343958 364350
rect 343338 364226 343958 364294
rect 343338 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 343958 364226
rect 343338 364102 343958 364170
rect 343338 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 343958 364102
rect 343338 363978 343958 364046
rect 343338 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 343958 363978
rect 343338 346350 343958 363922
rect 343338 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 343958 346350
rect 343338 346226 343958 346294
rect 343338 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 343958 346226
rect 343338 346102 343958 346170
rect 343338 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 343958 346102
rect 343338 345978 343958 346046
rect 343338 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 343958 345978
rect 343338 328350 343958 345922
rect 343338 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 343958 328350
rect 343338 328226 343958 328294
rect 343338 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 343958 328226
rect 343338 328102 343958 328170
rect 343338 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 343958 328102
rect 343338 327978 343958 328046
rect 343338 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 343958 327978
rect 343338 310350 343958 327922
rect 343338 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 343958 310350
rect 343338 310226 343958 310294
rect 343338 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 343958 310226
rect 343338 310102 343958 310170
rect 343338 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 343958 310102
rect 343338 309978 343958 310046
rect 343338 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 343958 309978
rect 343338 292350 343958 309922
rect 343338 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 343958 292350
rect 343338 292226 343958 292294
rect 343338 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 343958 292226
rect 343338 292102 343958 292170
rect 343338 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 343958 292102
rect 343338 291978 343958 292046
rect 343338 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 343958 291978
rect 343338 274350 343958 291922
rect 343338 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 343958 274350
rect 343338 274226 343958 274294
rect 343338 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 343958 274226
rect 343338 274102 343958 274170
rect 343338 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 343958 274102
rect 343338 273978 343958 274046
rect 343338 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 343958 273978
rect 343338 256350 343958 273922
rect 343338 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 343958 256350
rect 343338 256226 343958 256294
rect 343338 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 343958 256226
rect 343338 256102 343958 256170
rect 343338 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 343958 256102
rect 343338 255978 343958 256046
rect 343338 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 343958 255978
rect 343338 238350 343958 255922
rect 343338 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 343958 238350
rect 343338 238226 343958 238294
rect 343338 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 343958 238226
rect 343338 238102 343958 238170
rect 343338 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 343958 238102
rect 343338 237978 343958 238046
rect 343338 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 343958 237978
rect 343338 220350 343958 237922
rect 343338 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 343958 220350
rect 343338 220226 343958 220294
rect 343338 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 343958 220226
rect 343338 220102 343958 220170
rect 343338 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 343958 220102
rect 343338 219978 343958 220046
rect 343338 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 343958 219978
rect 343338 202350 343958 219922
rect 343338 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 343958 202350
rect 343338 202226 343958 202294
rect 343338 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 343958 202226
rect 343338 202102 343958 202170
rect 343338 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 343958 202102
rect 343338 201978 343958 202046
rect 343338 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 343958 201978
rect 343338 184350 343958 201922
rect 343338 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 343958 184350
rect 343338 184226 343958 184294
rect 343338 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 343958 184226
rect 343338 184102 343958 184170
rect 343338 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 343958 184102
rect 343338 183978 343958 184046
rect 343338 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 343958 183978
rect 343338 166350 343958 183922
rect 343338 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 343958 166350
rect 343338 166226 343958 166294
rect 343338 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 343958 166226
rect 343338 166102 343958 166170
rect 343338 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 343958 166102
rect 343338 165978 343958 166046
rect 343338 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 343958 165978
rect 329308 163828 329364 163838
rect 316338 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 316958 154350
rect 316338 154226 316958 154294
rect 316338 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 316958 154226
rect 316338 154102 316958 154170
rect 316338 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 316958 154102
rect 316338 153978 316958 154046
rect 316338 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 316958 153978
rect 314636 141204 314692 141214
rect 314636 141058 314692 141148
rect 314636 140992 314692 141002
rect 312618 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 313238 130350
rect 312618 130226 313238 130294
rect 312618 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 313238 130226
rect 312618 130102 313238 130170
rect 312618 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 313238 130102
rect 312618 129978 313238 130046
rect 312618 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 313238 129978
rect 312618 112350 313238 129922
rect 312618 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 313238 112350
rect 312618 112226 313238 112294
rect 312618 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 313238 112226
rect 312618 112102 313238 112170
rect 312618 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 313238 112102
rect 312618 111978 313238 112046
rect 312618 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 313238 111978
rect 312618 94350 313238 111922
rect 312618 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 313238 94350
rect 312618 94226 313238 94294
rect 312618 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 313238 94226
rect 312618 94102 313238 94170
rect 312618 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 313238 94102
rect 312618 93978 313238 94046
rect 312618 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 313238 93978
rect 312618 76350 313238 93922
rect 312618 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 313238 76350
rect 312618 76226 313238 76294
rect 312618 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 313238 76226
rect 312618 76102 313238 76170
rect 312618 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 313238 76102
rect 312618 75978 313238 76046
rect 312618 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 313238 75978
rect 312618 58350 313238 75922
rect 312618 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 313238 58350
rect 312618 58226 313238 58294
rect 312618 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 313238 58226
rect 312618 58102 313238 58170
rect 312618 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 313238 58102
rect 312618 57978 313238 58046
rect 312618 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 313238 57978
rect 312618 40350 313238 57922
rect 312618 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 313238 40350
rect 312618 40226 313238 40294
rect 312618 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 313238 40226
rect 312618 40102 313238 40170
rect 312618 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 313238 40102
rect 312618 39978 313238 40046
rect 312618 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 313238 39978
rect 312618 22350 313238 39922
rect 312618 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 313238 22350
rect 312618 22226 313238 22294
rect 312618 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 313238 22226
rect 312618 22102 313238 22170
rect 312618 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 313238 22102
rect 312618 21978 313238 22046
rect 312618 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 313238 21978
rect 312618 4350 313238 21922
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 285618 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 286238 -1120
rect 285618 -1244 286238 -1176
rect 285618 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 286238 -1244
rect 285618 -1368 286238 -1300
rect 285618 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 286238 -1368
rect 285618 -1492 286238 -1424
rect 285618 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 286238 -1492
rect 285618 -1644 286238 -1548
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 316338 136350 316958 153922
rect 322588 162148 322644 162158
rect 319228 141958 319284 141968
rect 319228 141204 319284 141902
rect 319228 141138 319284 141148
rect 316338 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 316958 136350
rect 316338 136226 316958 136294
rect 316338 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 316958 136226
rect 316338 136102 316958 136170
rect 316338 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 316958 136102
rect 316338 135978 316958 136046
rect 316338 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 316958 135978
rect 316338 118350 316958 135922
rect 316338 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 316958 118350
rect 316338 118226 316958 118294
rect 316338 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 316958 118226
rect 316338 118102 316958 118170
rect 316338 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 316958 118102
rect 316338 117978 316958 118046
rect 316338 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 316958 117978
rect 316338 100350 316958 117922
rect 316338 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 316958 100350
rect 316338 100226 316958 100294
rect 316338 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 316958 100226
rect 316338 100102 316958 100170
rect 316338 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 316958 100102
rect 316338 99978 316958 100046
rect 316338 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 316958 99978
rect 316338 82350 316958 99922
rect 316338 82294 316434 82350
rect 316490 82294 316558 82350
rect 316614 82294 316682 82350
rect 316738 82294 316806 82350
rect 316862 82294 316958 82350
rect 316338 82226 316958 82294
rect 316338 82170 316434 82226
rect 316490 82170 316558 82226
rect 316614 82170 316682 82226
rect 316738 82170 316806 82226
rect 316862 82170 316958 82226
rect 316338 82102 316958 82170
rect 316338 82046 316434 82102
rect 316490 82046 316558 82102
rect 316614 82046 316682 82102
rect 316738 82046 316806 82102
rect 316862 82046 316958 82102
rect 316338 81978 316958 82046
rect 316338 81922 316434 81978
rect 316490 81922 316558 81978
rect 316614 81922 316682 81978
rect 316738 81922 316806 81978
rect 316862 81922 316958 81978
rect 316338 64350 316958 81922
rect 316338 64294 316434 64350
rect 316490 64294 316558 64350
rect 316614 64294 316682 64350
rect 316738 64294 316806 64350
rect 316862 64294 316958 64350
rect 316338 64226 316958 64294
rect 316338 64170 316434 64226
rect 316490 64170 316558 64226
rect 316614 64170 316682 64226
rect 316738 64170 316806 64226
rect 316862 64170 316958 64226
rect 316338 64102 316958 64170
rect 316338 64046 316434 64102
rect 316490 64046 316558 64102
rect 316614 64046 316682 64102
rect 316738 64046 316806 64102
rect 316862 64046 316958 64102
rect 316338 63978 316958 64046
rect 316338 63922 316434 63978
rect 316490 63922 316558 63978
rect 316614 63922 316682 63978
rect 316738 63922 316806 63978
rect 316862 63922 316958 63978
rect 316338 46350 316958 63922
rect 316338 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 316958 46350
rect 316338 46226 316958 46294
rect 316338 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 316958 46226
rect 316338 46102 316958 46170
rect 316338 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 316958 46102
rect 316338 45978 316958 46046
rect 316338 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 316958 45978
rect 316338 28350 316958 45922
rect 316338 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 316958 28350
rect 316338 28226 316958 28294
rect 316338 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 316958 28226
rect 316338 28102 316958 28170
rect 316338 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 316958 28102
rect 316338 27978 316958 28046
rect 316338 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 316958 27978
rect 316338 10350 316958 27922
rect 316338 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 316958 10350
rect 316338 10226 316958 10294
rect 316338 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 316958 10226
rect 316338 10102 316958 10170
rect 316338 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 316958 10102
rect 316338 9978 316958 10046
rect 316338 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 316958 9978
rect 316338 -1120 316958 9922
rect 322588 4228 322644 162092
rect 322588 4162 322644 4172
rect 329308 4228 329364 163772
rect 343338 148350 343958 165922
rect 343338 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 343958 148350
rect 343338 148226 343958 148294
rect 343338 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 343958 148226
rect 343338 148102 343958 148170
rect 343338 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 343958 148102
rect 343338 147978 343958 148046
rect 343338 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 343958 147978
rect 330876 142772 330932 142782
rect 330876 141958 330932 142716
rect 330876 141892 330932 141902
rect 333452 142772 333508 142782
rect 333452 141058 333508 142716
rect 333452 140992 333508 141002
rect 340956 141204 341012 141214
rect 340956 140878 341012 141148
rect 340956 140812 341012 140822
rect 329308 4162 329364 4172
rect 343338 130350 343958 147922
rect 347058 388350 347678 402722
rect 347058 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 347678 388350
rect 347058 388226 347678 388294
rect 347058 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 347678 388226
rect 347058 388102 347678 388170
rect 347058 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 347678 388102
rect 347058 387978 347678 388046
rect 347058 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 347678 387978
rect 347058 370350 347678 387922
rect 347058 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 347678 370350
rect 347058 370226 347678 370294
rect 347058 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 347678 370226
rect 347058 370102 347678 370170
rect 347058 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 347678 370102
rect 347058 369978 347678 370046
rect 347058 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 347678 369978
rect 347058 352350 347678 369922
rect 347058 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 347678 352350
rect 347058 352226 347678 352294
rect 347058 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 347678 352226
rect 347058 352102 347678 352170
rect 347058 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 347678 352102
rect 347058 351978 347678 352046
rect 347058 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 347678 351978
rect 347058 334350 347678 351922
rect 374058 400350 374678 402722
rect 374058 400294 374154 400350
rect 374210 400294 374278 400350
rect 374334 400294 374402 400350
rect 374458 400294 374526 400350
rect 374582 400294 374678 400350
rect 374058 400226 374678 400294
rect 374058 400170 374154 400226
rect 374210 400170 374278 400226
rect 374334 400170 374402 400226
rect 374458 400170 374526 400226
rect 374582 400170 374678 400226
rect 374058 400102 374678 400170
rect 374058 400046 374154 400102
rect 374210 400046 374278 400102
rect 374334 400046 374402 400102
rect 374458 400046 374526 400102
rect 374582 400046 374678 400102
rect 374058 399978 374678 400046
rect 374058 399922 374154 399978
rect 374210 399922 374278 399978
rect 374334 399922 374402 399978
rect 374458 399922 374526 399978
rect 374582 399922 374678 399978
rect 374058 382350 374678 399922
rect 374058 382294 374154 382350
rect 374210 382294 374278 382350
rect 374334 382294 374402 382350
rect 374458 382294 374526 382350
rect 374582 382294 374678 382350
rect 374058 382226 374678 382294
rect 374058 382170 374154 382226
rect 374210 382170 374278 382226
rect 374334 382170 374402 382226
rect 374458 382170 374526 382226
rect 374582 382170 374678 382226
rect 374058 382102 374678 382170
rect 374058 382046 374154 382102
rect 374210 382046 374278 382102
rect 374334 382046 374402 382102
rect 374458 382046 374526 382102
rect 374582 382046 374678 382102
rect 374058 381978 374678 382046
rect 374058 381922 374154 381978
rect 374210 381922 374278 381978
rect 374334 381922 374402 381978
rect 374458 381922 374526 381978
rect 374582 381922 374678 381978
rect 374058 364350 374678 381922
rect 374058 364294 374154 364350
rect 374210 364294 374278 364350
rect 374334 364294 374402 364350
rect 374458 364294 374526 364350
rect 374582 364294 374678 364350
rect 374058 364226 374678 364294
rect 374058 364170 374154 364226
rect 374210 364170 374278 364226
rect 374334 364170 374402 364226
rect 374458 364170 374526 364226
rect 374582 364170 374678 364226
rect 374058 364102 374678 364170
rect 374058 364046 374154 364102
rect 374210 364046 374278 364102
rect 374334 364046 374402 364102
rect 374458 364046 374526 364102
rect 374582 364046 374678 364102
rect 374058 363978 374678 364046
rect 374058 363922 374154 363978
rect 374210 363922 374278 363978
rect 374334 363922 374402 363978
rect 374458 363922 374526 363978
rect 374582 363922 374678 363978
rect 347058 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 347678 334350
rect 347058 334226 347678 334294
rect 347058 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 347678 334226
rect 347058 334102 347678 334170
rect 347058 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 347678 334102
rect 347058 333978 347678 334046
rect 347058 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 347678 333978
rect 347058 316350 347678 333922
rect 355292 349498 355348 349508
rect 351932 330058 351988 330068
rect 347058 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 347678 316350
rect 347058 316226 347678 316294
rect 347058 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 347678 316226
rect 347058 316102 347678 316170
rect 347058 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 347678 316102
rect 347058 315978 347678 316046
rect 347058 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 347678 315978
rect 347058 298350 347678 315922
rect 347058 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 347678 298350
rect 347058 298226 347678 298294
rect 347058 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 347678 298226
rect 347058 298102 347678 298170
rect 347058 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 347678 298102
rect 347058 297978 347678 298046
rect 347058 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 347678 297978
rect 347058 280350 347678 297922
rect 347058 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 347678 280350
rect 347058 280226 347678 280294
rect 347058 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 347678 280226
rect 347058 280102 347678 280170
rect 347058 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 347678 280102
rect 347058 279978 347678 280046
rect 347058 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 347678 279978
rect 347058 262350 347678 279922
rect 347058 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 347678 262350
rect 347058 262226 347678 262294
rect 347058 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 347678 262226
rect 347058 262102 347678 262170
rect 347058 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 347678 262102
rect 347058 261978 347678 262046
rect 347058 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 347678 261978
rect 347058 244350 347678 261922
rect 347058 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 347678 244350
rect 347058 244226 347678 244294
rect 347058 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 347678 244226
rect 347058 244102 347678 244170
rect 347058 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 347678 244102
rect 347058 243978 347678 244046
rect 347058 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 347678 243978
rect 347058 226350 347678 243922
rect 347058 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 347678 226350
rect 347058 226226 347678 226294
rect 347058 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 347678 226226
rect 347058 226102 347678 226170
rect 347058 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 347678 226102
rect 347058 225978 347678 226046
rect 347058 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 347678 225978
rect 347058 208350 347678 225922
rect 347058 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 347678 208350
rect 347058 208226 347678 208294
rect 347058 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 347678 208226
rect 347058 208102 347678 208170
rect 347058 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 347678 208102
rect 347058 207978 347678 208046
rect 347058 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 347678 207978
rect 347058 190350 347678 207922
rect 347058 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 347678 190350
rect 347058 190226 347678 190294
rect 347058 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 347678 190226
rect 347058 190102 347678 190170
rect 347058 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 347678 190102
rect 347058 189978 347678 190046
rect 347058 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 347678 189978
rect 347058 172350 347678 189922
rect 347058 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 347678 172350
rect 347058 172226 347678 172294
rect 347058 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 347678 172226
rect 347058 172102 347678 172170
rect 347058 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 347678 172102
rect 347058 171978 347678 172046
rect 347058 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 347678 171978
rect 347058 154350 347678 171922
rect 347058 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 347678 154350
rect 347058 154226 347678 154294
rect 347058 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 347678 154226
rect 347058 154102 347678 154170
rect 347058 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 347678 154102
rect 347058 153978 347678 154046
rect 347058 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 347678 153978
rect 344652 142138 344708 142148
rect 344652 142034 344708 142044
rect 347058 137760 347678 153922
rect 348572 319978 348628 319988
rect 343338 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 343958 130350
rect 343338 130226 343958 130294
rect 343338 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 343958 130226
rect 343338 130102 343958 130170
rect 343338 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 343958 130102
rect 343338 129978 343958 130046
rect 343338 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 343958 129978
rect 343338 112350 343958 129922
rect 345788 130350 346264 130384
rect 345788 130294 345812 130350
rect 345868 130294 345936 130350
rect 345992 130294 346060 130350
rect 346116 130294 346184 130350
rect 346240 130294 346264 130350
rect 345788 130226 346264 130294
rect 345788 130170 345812 130226
rect 345868 130170 345936 130226
rect 345992 130170 346060 130226
rect 346116 130170 346184 130226
rect 346240 130170 346264 130226
rect 345788 130102 346264 130170
rect 345788 130046 345812 130102
rect 345868 130046 345936 130102
rect 345992 130046 346060 130102
rect 346116 130046 346184 130102
rect 346240 130046 346264 130102
rect 345788 129978 346264 130046
rect 345788 129922 345812 129978
rect 345868 129922 345936 129978
rect 345992 129922 346060 129978
rect 346116 129922 346184 129978
rect 346240 129922 346264 129978
rect 345788 129888 346264 129922
rect 346588 118350 347064 118384
rect 346588 118294 346612 118350
rect 346668 118294 346736 118350
rect 346792 118294 346860 118350
rect 346916 118294 346984 118350
rect 347040 118294 347064 118350
rect 346588 118226 347064 118294
rect 346588 118170 346612 118226
rect 346668 118170 346736 118226
rect 346792 118170 346860 118226
rect 346916 118170 346984 118226
rect 347040 118170 347064 118226
rect 346588 118102 347064 118170
rect 346588 118046 346612 118102
rect 346668 118046 346736 118102
rect 346792 118046 346860 118102
rect 346916 118046 346984 118102
rect 347040 118046 347064 118102
rect 346588 117978 347064 118046
rect 346588 117922 346612 117978
rect 346668 117922 346736 117978
rect 346792 117922 346860 117978
rect 346916 117922 346984 117978
rect 347040 117922 347064 117978
rect 346588 117888 347064 117922
rect 343338 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 343958 112350
rect 343338 112226 343958 112294
rect 343338 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 343958 112226
rect 343338 112102 343958 112170
rect 343338 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 343958 112102
rect 343338 111978 343958 112046
rect 343338 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 343958 111978
rect 343338 94350 343958 111922
rect 345788 112350 346264 112384
rect 345788 112294 345812 112350
rect 345868 112294 345936 112350
rect 345992 112294 346060 112350
rect 346116 112294 346184 112350
rect 346240 112294 346264 112350
rect 345788 112226 346264 112294
rect 345788 112170 345812 112226
rect 345868 112170 345936 112226
rect 345992 112170 346060 112226
rect 346116 112170 346184 112226
rect 346240 112170 346264 112226
rect 345788 112102 346264 112170
rect 345788 112046 345812 112102
rect 345868 112046 345936 112102
rect 345992 112046 346060 112102
rect 346116 112046 346184 112102
rect 346240 112046 346264 112102
rect 345788 111978 346264 112046
rect 345788 111922 345812 111978
rect 345868 111922 345936 111978
rect 345992 111922 346060 111978
rect 346116 111922 346184 111978
rect 346240 111922 346264 111978
rect 345788 111888 346264 111922
rect 346588 100350 347064 100384
rect 346588 100294 346612 100350
rect 346668 100294 346736 100350
rect 346792 100294 346860 100350
rect 346916 100294 346984 100350
rect 347040 100294 347064 100350
rect 346588 100226 347064 100294
rect 346588 100170 346612 100226
rect 346668 100170 346736 100226
rect 346792 100170 346860 100226
rect 346916 100170 346984 100226
rect 347040 100170 347064 100226
rect 346588 100102 347064 100170
rect 346588 100046 346612 100102
rect 346668 100046 346736 100102
rect 346792 100046 346860 100102
rect 346916 100046 346984 100102
rect 347040 100046 347064 100102
rect 346588 99978 347064 100046
rect 346588 99922 346612 99978
rect 346668 99922 346736 99978
rect 346792 99922 346860 99978
rect 346916 99922 346984 99978
rect 347040 99922 347064 99978
rect 346588 99888 347064 99922
rect 343338 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 343958 94350
rect 343338 94226 343958 94294
rect 343338 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 343958 94226
rect 343338 94102 343958 94170
rect 343338 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 343958 94102
rect 343338 93978 343958 94046
rect 343338 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 343958 93978
rect 343338 76350 343958 93922
rect 345788 94350 346264 94384
rect 345788 94294 345812 94350
rect 345868 94294 345936 94350
rect 345992 94294 346060 94350
rect 346116 94294 346184 94350
rect 346240 94294 346264 94350
rect 345788 94226 346264 94294
rect 345788 94170 345812 94226
rect 345868 94170 345936 94226
rect 345992 94170 346060 94226
rect 346116 94170 346184 94226
rect 346240 94170 346264 94226
rect 345788 94102 346264 94170
rect 345788 94046 345812 94102
rect 345868 94046 345936 94102
rect 345992 94046 346060 94102
rect 346116 94046 346184 94102
rect 346240 94046 346264 94102
rect 345788 93978 346264 94046
rect 345788 93922 345812 93978
rect 345868 93922 345936 93978
rect 345992 93922 346060 93978
rect 346116 93922 346184 93978
rect 346240 93922 346264 93978
rect 345788 93888 346264 93922
rect 346588 82350 347064 82384
rect 346588 82294 346612 82350
rect 346668 82294 346736 82350
rect 346792 82294 346860 82350
rect 346916 82294 346984 82350
rect 347040 82294 347064 82350
rect 346588 82226 347064 82294
rect 346588 82170 346612 82226
rect 346668 82170 346736 82226
rect 346792 82170 346860 82226
rect 346916 82170 346984 82226
rect 347040 82170 347064 82226
rect 346588 82102 347064 82170
rect 346588 82046 346612 82102
rect 346668 82046 346736 82102
rect 346792 82046 346860 82102
rect 346916 82046 346984 82102
rect 347040 82046 347064 82102
rect 346588 81978 347064 82046
rect 346588 81922 346612 81978
rect 346668 81922 346736 81978
rect 346792 81922 346860 81978
rect 346916 81922 346984 81978
rect 347040 81922 347064 81978
rect 346588 81888 347064 81922
rect 343338 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 343958 76350
rect 343338 76226 343958 76294
rect 343338 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 343958 76226
rect 343338 76102 343958 76170
rect 343338 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 343958 76102
rect 343338 75978 343958 76046
rect 343338 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 343958 75978
rect 343338 58350 343958 75922
rect 345788 76350 346264 76384
rect 345788 76294 345812 76350
rect 345868 76294 345936 76350
rect 345992 76294 346060 76350
rect 346116 76294 346184 76350
rect 346240 76294 346264 76350
rect 345788 76226 346264 76294
rect 345788 76170 345812 76226
rect 345868 76170 345936 76226
rect 345992 76170 346060 76226
rect 346116 76170 346184 76226
rect 346240 76170 346264 76226
rect 345788 76102 346264 76170
rect 345788 76046 345812 76102
rect 345868 76046 345936 76102
rect 345992 76046 346060 76102
rect 346116 76046 346184 76102
rect 346240 76046 346264 76102
rect 345788 75978 346264 76046
rect 345788 75922 345812 75978
rect 345868 75922 345936 75978
rect 345992 75922 346060 75978
rect 346116 75922 346184 75978
rect 346240 75922 346264 75978
rect 345788 75888 346264 75922
rect 346588 64350 347064 64384
rect 346588 64294 346612 64350
rect 346668 64294 346736 64350
rect 346792 64294 346860 64350
rect 346916 64294 346984 64350
rect 347040 64294 347064 64350
rect 346588 64226 347064 64294
rect 346588 64170 346612 64226
rect 346668 64170 346736 64226
rect 346792 64170 346860 64226
rect 346916 64170 346984 64226
rect 347040 64170 347064 64226
rect 346588 64102 347064 64170
rect 346588 64046 346612 64102
rect 346668 64046 346736 64102
rect 346792 64046 346860 64102
rect 346916 64046 346984 64102
rect 347040 64046 347064 64102
rect 346588 63978 347064 64046
rect 346588 63922 346612 63978
rect 346668 63922 346736 63978
rect 346792 63922 346860 63978
rect 346916 63922 346984 63978
rect 347040 63922 347064 63978
rect 346588 63888 347064 63922
rect 343338 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 343958 58350
rect 343338 58226 343958 58294
rect 343338 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 343958 58226
rect 343338 58102 343958 58170
rect 343338 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 343958 58102
rect 343338 57978 343958 58046
rect 343338 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 343958 57978
rect 343338 40350 343958 57922
rect 345788 58350 346264 58384
rect 345788 58294 345812 58350
rect 345868 58294 345936 58350
rect 345992 58294 346060 58350
rect 346116 58294 346184 58350
rect 346240 58294 346264 58350
rect 345788 58226 346264 58294
rect 345788 58170 345812 58226
rect 345868 58170 345936 58226
rect 345992 58170 346060 58226
rect 346116 58170 346184 58226
rect 346240 58170 346264 58226
rect 345788 58102 346264 58170
rect 345788 58046 345812 58102
rect 345868 58046 345936 58102
rect 345992 58046 346060 58102
rect 346116 58046 346184 58102
rect 346240 58046 346264 58102
rect 345788 57978 346264 58046
rect 345788 57922 345812 57978
rect 345868 57922 345936 57978
rect 345992 57922 346060 57978
rect 346116 57922 346184 57978
rect 346240 57922 346264 57978
rect 345788 57888 346264 57922
rect 346588 46350 347064 46384
rect 346588 46294 346612 46350
rect 346668 46294 346736 46350
rect 346792 46294 346860 46350
rect 346916 46294 346984 46350
rect 347040 46294 347064 46350
rect 346588 46226 347064 46294
rect 346588 46170 346612 46226
rect 346668 46170 346736 46226
rect 346792 46170 346860 46226
rect 346916 46170 346984 46226
rect 347040 46170 347064 46226
rect 346588 46102 347064 46170
rect 346588 46046 346612 46102
rect 346668 46046 346736 46102
rect 346792 46046 346860 46102
rect 346916 46046 346984 46102
rect 347040 46046 347064 46102
rect 346588 45978 347064 46046
rect 346588 45922 346612 45978
rect 346668 45922 346736 45978
rect 346792 45922 346860 45978
rect 346916 45922 346984 45978
rect 347040 45922 347064 45978
rect 346588 45888 347064 45922
rect 343338 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 343958 40350
rect 343338 40226 343958 40294
rect 343338 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 343958 40226
rect 343338 40102 343958 40170
rect 343338 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 343958 40102
rect 343338 39978 343958 40046
rect 343338 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 343958 39978
rect 343338 22350 343958 39922
rect 343338 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 343958 22350
rect 343338 22226 343958 22294
rect 343338 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 343958 22226
rect 343338 22102 343958 22170
rect 343338 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 343958 22102
rect 343338 21978 343958 22046
rect 343338 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 343958 21978
rect 343338 4350 343958 21922
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 316338 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 316958 -1120
rect 316338 -1244 316958 -1176
rect 316338 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 316958 -1244
rect 316338 -1368 316958 -1300
rect 316338 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 316958 -1368
rect 316338 -1492 316958 -1424
rect 316338 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 316958 -1492
rect 316338 -1644 316958 -1548
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 347058 28350 347678 41024
rect 347058 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 347678 28350
rect 347058 28226 347678 28294
rect 347058 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 347678 28226
rect 347058 28102 347678 28170
rect 347058 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 347678 28102
rect 347058 27978 347678 28046
rect 347058 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 347678 27978
rect 347058 10350 347678 27922
rect 347058 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 347678 10350
rect 347058 10226 347678 10294
rect 347058 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 347678 10226
rect 347058 10102 347678 10170
rect 347058 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 347678 10102
rect 347058 9978 347678 10046
rect 347058 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 347678 9978
rect 347058 -1120 347678 9922
rect 348572 4340 348628 319922
rect 350252 311698 350308 311708
rect 350252 4788 350308 311642
rect 350252 4722 350308 4732
rect 351932 4452 351988 330002
rect 353612 325018 353668 325028
rect 353612 4676 353668 324962
rect 355292 36148 355348 349442
rect 374058 346350 374678 363922
rect 374058 346294 374154 346350
rect 374210 346294 374278 346350
rect 374334 346294 374402 346350
rect 374458 346294 374526 346350
rect 374582 346294 374678 346350
rect 374058 346226 374678 346294
rect 374058 346170 374154 346226
rect 374210 346170 374278 346226
rect 374334 346170 374402 346226
rect 374458 346170 374526 346226
rect 374582 346170 374678 346226
rect 374058 346102 374678 346170
rect 374058 346046 374154 346102
rect 374210 346046 374278 346102
rect 374334 346046 374402 346102
rect 374458 346046 374526 346102
rect 374582 346046 374678 346102
rect 374058 345978 374678 346046
rect 374058 345922 374154 345978
rect 374210 345922 374278 345978
rect 374334 345922 374402 345978
rect 374458 345922 374526 345978
rect 374582 345922 374678 345978
rect 355292 36082 355348 36092
rect 358652 343738 358708 343748
rect 353612 4610 353668 4620
rect 351932 4386 351988 4396
rect 348572 4274 348628 4284
rect 358652 4228 358708 343682
rect 374058 328350 374678 345922
rect 374058 328294 374154 328350
rect 374210 328294 374278 328350
rect 374334 328294 374402 328350
rect 374458 328294 374526 328350
rect 374582 328294 374678 328350
rect 374058 328226 374678 328294
rect 374058 328170 374154 328226
rect 374210 328170 374278 328226
rect 374334 328170 374402 328226
rect 374458 328170 374526 328226
rect 374582 328170 374678 328226
rect 374058 328102 374678 328170
rect 374058 328046 374154 328102
rect 374210 328046 374278 328102
rect 374334 328046 374402 328102
rect 374458 328046 374526 328102
rect 374582 328046 374678 328102
rect 374058 327978 374678 328046
rect 374058 327922 374154 327978
rect 374210 327922 374278 327978
rect 374334 327922 374402 327978
rect 374458 327922 374526 327978
rect 374582 327922 374678 327978
rect 360332 323398 360388 323408
rect 360332 4564 360388 323342
rect 374058 310350 374678 327922
rect 374058 310294 374154 310350
rect 374210 310294 374278 310350
rect 374334 310294 374402 310350
rect 374458 310294 374526 310350
rect 374582 310294 374678 310350
rect 374058 310226 374678 310294
rect 374058 310170 374154 310226
rect 374210 310170 374278 310226
rect 374334 310170 374402 310226
rect 374458 310170 374526 310226
rect 374582 310170 374678 310226
rect 374058 310102 374678 310170
rect 374058 310046 374154 310102
rect 374210 310046 374278 310102
rect 374334 310046 374402 310102
rect 374458 310046 374526 310102
rect 374582 310046 374678 310102
rect 374058 309978 374678 310046
rect 374058 309922 374154 309978
rect 374210 309922 374278 309978
rect 374334 309922 374402 309978
rect 374458 309922 374526 309978
rect 374582 309922 374678 309978
rect 374058 292350 374678 309922
rect 374058 292294 374154 292350
rect 374210 292294 374278 292350
rect 374334 292294 374402 292350
rect 374458 292294 374526 292350
rect 374582 292294 374678 292350
rect 374058 292226 374678 292294
rect 374058 292170 374154 292226
rect 374210 292170 374278 292226
rect 374334 292170 374402 292226
rect 374458 292170 374526 292226
rect 374582 292170 374678 292226
rect 374058 292102 374678 292170
rect 374058 292046 374154 292102
rect 374210 292046 374278 292102
rect 374334 292046 374402 292102
rect 374458 292046 374526 292102
rect 374582 292046 374678 292102
rect 374058 291978 374678 292046
rect 374058 291922 374154 291978
rect 374210 291922 374278 291978
rect 374334 291922 374402 291978
rect 374458 291922 374526 291978
rect 374582 291922 374678 291978
rect 374058 274350 374678 291922
rect 374058 274294 374154 274350
rect 374210 274294 374278 274350
rect 374334 274294 374402 274350
rect 374458 274294 374526 274350
rect 374582 274294 374678 274350
rect 374058 274226 374678 274294
rect 374058 274170 374154 274226
rect 374210 274170 374278 274226
rect 374334 274170 374402 274226
rect 374458 274170 374526 274226
rect 374582 274170 374678 274226
rect 374058 274102 374678 274170
rect 374058 274046 374154 274102
rect 374210 274046 374278 274102
rect 374334 274046 374402 274102
rect 374458 274046 374526 274102
rect 374582 274046 374678 274102
rect 374058 273978 374678 274046
rect 374058 273922 374154 273978
rect 374210 273922 374278 273978
rect 374334 273922 374402 273978
rect 374458 273922 374526 273978
rect 374582 273922 374678 273978
rect 364252 259140 364308 259150
rect 363916 258692 363972 258702
rect 361906 244350 362382 244384
rect 361906 244294 361930 244350
rect 361986 244294 362054 244350
rect 362110 244294 362178 244350
rect 362234 244294 362302 244350
rect 362358 244294 362382 244350
rect 361906 244226 362382 244294
rect 361906 244170 361930 244226
rect 361986 244170 362054 244226
rect 362110 244170 362178 244226
rect 362234 244170 362302 244226
rect 362358 244170 362382 244226
rect 361906 244102 362382 244170
rect 361906 244046 361930 244102
rect 361986 244046 362054 244102
rect 362110 244046 362178 244102
rect 362234 244046 362302 244102
rect 362358 244046 362382 244102
rect 361906 243978 362382 244046
rect 361906 243922 361930 243978
rect 361986 243922 362054 243978
rect 362110 243922 362178 243978
rect 362234 243922 362302 243978
rect 362358 243922 362382 243978
rect 361906 243888 362382 243922
rect 363916 243628 363972 258636
rect 363692 243572 363972 243628
rect 361106 238350 361582 238384
rect 361106 238294 361130 238350
rect 361186 238294 361254 238350
rect 361310 238294 361378 238350
rect 361434 238294 361502 238350
rect 361558 238294 361582 238350
rect 361106 238226 361582 238294
rect 361106 238170 361130 238226
rect 361186 238170 361254 238226
rect 361310 238170 361378 238226
rect 361434 238170 361502 238226
rect 361558 238170 361582 238226
rect 361106 238102 361582 238170
rect 361106 238046 361130 238102
rect 361186 238046 361254 238102
rect 361310 238046 361378 238102
rect 361434 238046 361502 238102
rect 361558 238046 361582 238102
rect 361106 237978 361582 238046
rect 361106 237922 361130 237978
rect 361186 237922 361254 237978
rect 361310 237922 361378 237978
rect 361434 237922 361502 237978
rect 361558 237922 361582 237978
rect 361106 237888 361582 237922
rect 361906 226350 362382 226384
rect 361906 226294 361930 226350
rect 361986 226294 362054 226350
rect 362110 226294 362178 226350
rect 362234 226294 362302 226350
rect 362358 226294 362382 226350
rect 361906 226226 362382 226294
rect 361906 226170 361930 226226
rect 361986 226170 362054 226226
rect 362110 226170 362178 226226
rect 362234 226170 362302 226226
rect 362358 226170 362382 226226
rect 361906 226102 362382 226170
rect 361906 226046 361930 226102
rect 361986 226046 362054 226102
rect 362110 226046 362178 226102
rect 362234 226046 362302 226102
rect 362358 226046 362382 226102
rect 361906 225978 362382 226046
rect 361906 225922 361930 225978
rect 361986 225922 362054 225978
rect 362110 225922 362178 225978
rect 362234 225922 362302 225978
rect 362358 225922 362382 225978
rect 361906 225888 362382 225922
rect 361106 220350 361582 220384
rect 361106 220294 361130 220350
rect 361186 220294 361254 220350
rect 361310 220294 361378 220350
rect 361434 220294 361502 220350
rect 361558 220294 361582 220350
rect 361106 220226 361582 220294
rect 361106 220170 361130 220226
rect 361186 220170 361254 220226
rect 361310 220170 361378 220226
rect 361434 220170 361502 220226
rect 361558 220170 361582 220226
rect 361106 220102 361582 220170
rect 361106 220046 361130 220102
rect 361186 220046 361254 220102
rect 361310 220046 361378 220102
rect 361434 220046 361502 220102
rect 361558 220046 361582 220102
rect 361106 219978 361582 220046
rect 361106 219922 361130 219978
rect 361186 219922 361254 219978
rect 361310 219922 361378 219978
rect 361434 219922 361502 219978
rect 361558 219922 361582 219978
rect 361106 219888 361582 219922
rect 361906 208350 362382 208384
rect 361906 208294 361930 208350
rect 361986 208294 362054 208350
rect 362110 208294 362178 208350
rect 362234 208294 362302 208350
rect 362358 208294 362382 208350
rect 361906 208226 362382 208294
rect 361906 208170 361930 208226
rect 361986 208170 362054 208226
rect 362110 208170 362178 208226
rect 362234 208170 362302 208226
rect 362358 208170 362382 208226
rect 361906 208102 362382 208170
rect 361906 208046 361930 208102
rect 361986 208046 362054 208102
rect 362110 208046 362178 208102
rect 362234 208046 362302 208102
rect 362358 208046 362382 208102
rect 361906 207978 362382 208046
rect 361906 207922 361930 207978
rect 361986 207922 362054 207978
rect 362110 207922 362178 207978
rect 362234 207922 362302 207978
rect 362358 207922 362382 207978
rect 361906 207888 362382 207922
rect 361106 202350 361582 202384
rect 361106 202294 361130 202350
rect 361186 202294 361254 202350
rect 361310 202294 361378 202350
rect 361434 202294 361502 202350
rect 361558 202294 361582 202350
rect 361106 202226 361582 202294
rect 361106 202170 361130 202226
rect 361186 202170 361254 202226
rect 361310 202170 361378 202226
rect 361434 202170 361502 202226
rect 361558 202170 361582 202226
rect 361106 202102 361582 202170
rect 361106 202046 361130 202102
rect 361186 202046 361254 202102
rect 361310 202046 361378 202102
rect 361434 202046 361502 202102
rect 361558 202046 361582 202102
rect 361106 201978 361582 202046
rect 361106 201922 361130 201978
rect 361186 201922 361254 201978
rect 361310 201922 361378 201978
rect 361434 201922 361502 201978
rect 361558 201922 361582 201978
rect 361106 201888 361582 201922
rect 361906 190350 362382 190384
rect 361906 190294 361930 190350
rect 361986 190294 362054 190350
rect 362110 190294 362178 190350
rect 362234 190294 362302 190350
rect 362358 190294 362382 190350
rect 361906 190226 362382 190294
rect 361906 190170 361930 190226
rect 361986 190170 362054 190226
rect 362110 190170 362178 190226
rect 362234 190170 362302 190226
rect 362358 190170 362382 190226
rect 361906 190102 362382 190170
rect 361906 190046 361930 190102
rect 361986 190046 362054 190102
rect 362110 190046 362178 190102
rect 362234 190046 362302 190102
rect 362358 190046 362382 190102
rect 361906 189978 362382 190046
rect 361906 189922 361930 189978
rect 361986 189922 362054 189978
rect 362110 189922 362178 189978
rect 362234 189922 362302 189978
rect 362358 189922 362382 189978
rect 361906 189888 362382 189922
rect 361106 184350 361582 184384
rect 361106 184294 361130 184350
rect 361186 184294 361254 184350
rect 361310 184294 361378 184350
rect 361434 184294 361502 184350
rect 361558 184294 361582 184350
rect 361106 184226 361582 184294
rect 361106 184170 361130 184226
rect 361186 184170 361254 184226
rect 361310 184170 361378 184226
rect 361434 184170 361502 184226
rect 361558 184170 361582 184226
rect 361106 184102 361582 184170
rect 361106 184046 361130 184102
rect 361186 184046 361254 184102
rect 361310 184046 361378 184102
rect 361434 184046 361502 184102
rect 361558 184046 361582 184102
rect 361106 183978 361582 184046
rect 361106 183922 361130 183978
rect 361186 183922 361254 183978
rect 361310 183922 361378 183978
rect 361434 183922 361502 183978
rect 361558 183922 361582 183978
rect 361106 183888 361582 183922
rect 361906 172350 362382 172384
rect 361906 172294 361930 172350
rect 361986 172294 362054 172350
rect 362110 172294 362178 172350
rect 362234 172294 362302 172350
rect 362358 172294 362382 172350
rect 361906 172226 362382 172294
rect 361906 172170 361930 172226
rect 361986 172170 362054 172226
rect 362110 172170 362178 172226
rect 362234 172170 362302 172226
rect 362358 172170 362382 172226
rect 361906 172102 362382 172170
rect 361906 172046 361930 172102
rect 361986 172046 362054 172102
rect 362110 172046 362178 172102
rect 362234 172046 362302 172102
rect 362358 172046 362382 172102
rect 361906 171978 362382 172046
rect 361906 171922 361930 171978
rect 361986 171922 362054 171978
rect 362110 171922 362178 171978
rect 362234 171922 362302 171978
rect 362358 171922 362382 171978
rect 361906 171888 362382 171922
rect 361106 166350 361582 166384
rect 361106 166294 361130 166350
rect 361186 166294 361254 166350
rect 361310 166294 361378 166350
rect 361434 166294 361502 166350
rect 361558 166294 361582 166350
rect 361106 166226 361582 166294
rect 361106 166170 361130 166226
rect 361186 166170 361254 166226
rect 361310 166170 361378 166226
rect 361434 166170 361502 166226
rect 361558 166170 361582 166226
rect 361106 166102 361582 166170
rect 361106 166046 361130 166102
rect 361186 166046 361254 166102
rect 361310 166046 361378 166102
rect 361434 166046 361502 166102
rect 361558 166046 361582 166102
rect 361106 165978 361582 166046
rect 361106 165922 361130 165978
rect 361186 165922 361254 165978
rect 361310 165922 361378 165978
rect 361434 165922 361502 165978
rect 361558 165922 361582 165978
rect 361106 165888 361582 165922
rect 363692 141876 363748 243572
rect 364252 142324 364308 259084
rect 373884 259028 373940 259038
rect 373772 258692 373828 258702
rect 373772 149548 373828 258636
rect 364252 142258 364308 142268
rect 373436 149492 373828 149548
rect 363692 141810 363748 141820
rect 373436 141652 373492 149492
rect 373436 141204 373492 141596
rect 373436 141138 373492 141148
rect 373884 141092 373940 258972
rect 373884 139748 373940 141036
rect 373884 139682 373940 139692
rect 374058 256350 374678 273922
rect 377778 388350 378398 402722
rect 377778 388294 377874 388350
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 378398 388350
rect 377778 388226 378398 388294
rect 377778 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 378398 388226
rect 377778 388102 378398 388170
rect 377778 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 378398 388102
rect 377778 387978 378398 388046
rect 377778 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 378398 387978
rect 377778 370350 378398 387922
rect 404778 400350 405398 402722
rect 404778 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 405398 400350
rect 404778 400226 405398 400294
rect 404778 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 405398 400226
rect 404778 400102 405398 400170
rect 404778 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 405398 400102
rect 404778 399978 405398 400046
rect 404778 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 405398 399978
rect 404778 382350 405398 399922
rect 404778 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 405398 382350
rect 404778 382226 405398 382294
rect 404778 382170 404874 382226
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 405398 382226
rect 404778 382102 405398 382170
rect 404778 382046 404874 382102
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 405398 382102
rect 404778 381978 405398 382046
rect 404778 381922 404874 381978
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 405398 381978
rect 377778 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 378398 370350
rect 377778 370226 378398 370294
rect 377778 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 378398 370226
rect 377778 370102 378398 370170
rect 377778 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 378398 370102
rect 377778 369978 378398 370046
rect 377778 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 378398 369978
rect 377778 352350 378398 369922
rect 386590 370350 387066 370384
rect 386590 370294 386614 370350
rect 386670 370294 386738 370350
rect 386794 370294 386862 370350
rect 386918 370294 386986 370350
rect 387042 370294 387066 370350
rect 386590 370226 387066 370294
rect 386590 370170 386614 370226
rect 386670 370170 386738 370226
rect 386794 370170 386862 370226
rect 386918 370170 386986 370226
rect 387042 370170 387066 370226
rect 386590 370102 387066 370170
rect 386590 370046 386614 370102
rect 386670 370046 386738 370102
rect 386794 370046 386862 370102
rect 386918 370046 386986 370102
rect 387042 370046 387066 370102
rect 386590 369978 387066 370046
rect 386590 369922 386614 369978
rect 386670 369922 386738 369978
rect 386794 369922 386862 369978
rect 386918 369922 386986 369978
rect 387042 369922 387066 369978
rect 386590 369888 387066 369922
rect 387390 364350 387866 364384
rect 387390 364294 387414 364350
rect 387470 364294 387538 364350
rect 387594 364294 387662 364350
rect 387718 364294 387786 364350
rect 387842 364294 387866 364350
rect 387390 364226 387866 364294
rect 387390 364170 387414 364226
rect 387470 364170 387538 364226
rect 387594 364170 387662 364226
rect 387718 364170 387786 364226
rect 387842 364170 387866 364226
rect 387390 364102 387866 364170
rect 387390 364046 387414 364102
rect 387470 364046 387538 364102
rect 387594 364046 387662 364102
rect 387718 364046 387786 364102
rect 387842 364046 387866 364102
rect 387390 363978 387866 364046
rect 387390 363922 387414 363978
rect 387470 363922 387538 363978
rect 387594 363922 387662 363978
rect 387718 363922 387786 363978
rect 387842 363922 387866 363978
rect 387390 363888 387866 363922
rect 404778 364350 405398 381922
rect 404778 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 405398 364350
rect 404778 364226 405398 364294
rect 404778 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 405398 364226
rect 404778 364102 405398 364170
rect 404778 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 405398 364102
rect 404778 363978 405398 364046
rect 404778 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 405398 363978
rect 377778 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 378398 352350
rect 377778 352226 378398 352294
rect 377778 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 378398 352226
rect 377778 352102 378398 352170
rect 377778 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 378398 352102
rect 377778 351978 378398 352046
rect 377778 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 378398 351978
rect 377778 334350 378398 351922
rect 386590 352350 387066 352384
rect 386590 352294 386614 352350
rect 386670 352294 386738 352350
rect 386794 352294 386862 352350
rect 386918 352294 386986 352350
rect 387042 352294 387066 352350
rect 386590 352226 387066 352294
rect 386590 352170 386614 352226
rect 386670 352170 386738 352226
rect 386794 352170 386862 352226
rect 386918 352170 386986 352226
rect 387042 352170 387066 352226
rect 386590 352102 387066 352170
rect 386590 352046 386614 352102
rect 386670 352046 386738 352102
rect 386794 352046 386862 352102
rect 386918 352046 386986 352102
rect 387042 352046 387066 352102
rect 386590 351978 387066 352046
rect 386590 351922 386614 351978
rect 386670 351922 386738 351978
rect 386794 351922 386862 351978
rect 386918 351922 386986 351978
rect 387042 351922 387066 351978
rect 386590 351888 387066 351922
rect 387390 346350 387866 346384
rect 387390 346294 387414 346350
rect 387470 346294 387538 346350
rect 387594 346294 387662 346350
rect 387718 346294 387786 346350
rect 387842 346294 387866 346350
rect 387390 346226 387866 346294
rect 387390 346170 387414 346226
rect 387470 346170 387538 346226
rect 387594 346170 387662 346226
rect 387718 346170 387786 346226
rect 387842 346170 387866 346226
rect 387390 346102 387866 346170
rect 387390 346046 387414 346102
rect 387470 346046 387538 346102
rect 387594 346046 387662 346102
rect 387718 346046 387786 346102
rect 387842 346046 387866 346102
rect 387390 345978 387866 346046
rect 387390 345922 387414 345978
rect 387470 345922 387538 345978
rect 387594 345922 387662 345978
rect 387718 345922 387786 345978
rect 387842 345922 387866 345978
rect 387390 345888 387866 345922
rect 404778 346350 405398 363922
rect 404778 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 405398 346350
rect 404778 346226 405398 346294
rect 404778 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 405398 346226
rect 404778 346102 405398 346170
rect 404778 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 405398 346102
rect 404778 345978 405398 346046
rect 404778 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 405398 345978
rect 377778 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 378398 334350
rect 377778 334226 378398 334294
rect 377778 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 378398 334226
rect 377778 334102 378398 334170
rect 377778 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 378398 334102
rect 377778 333978 378398 334046
rect 377778 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 378398 333978
rect 377778 316350 378398 333922
rect 386590 334350 387066 334384
rect 386590 334294 386614 334350
rect 386670 334294 386738 334350
rect 386794 334294 386862 334350
rect 386918 334294 386986 334350
rect 387042 334294 387066 334350
rect 386590 334226 387066 334294
rect 386590 334170 386614 334226
rect 386670 334170 386738 334226
rect 386794 334170 386862 334226
rect 386918 334170 386986 334226
rect 387042 334170 387066 334226
rect 386590 334102 387066 334170
rect 386590 334046 386614 334102
rect 386670 334046 386738 334102
rect 386794 334046 386862 334102
rect 386918 334046 386986 334102
rect 387042 334046 387066 334102
rect 386590 333978 387066 334046
rect 386590 333922 386614 333978
rect 386670 333922 386738 333978
rect 386794 333922 386862 333978
rect 386918 333922 386986 333978
rect 387042 333922 387066 333978
rect 386590 333888 387066 333922
rect 390572 328580 390628 328590
rect 387390 328350 387866 328384
rect 387390 328294 387414 328350
rect 387470 328294 387538 328350
rect 387594 328294 387662 328350
rect 387718 328294 387786 328350
rect 387842 328294 387866 328350
rect 387390 328226 387866 328294
rect 387390 328170 387414 328226
rect 387470 328170 387538 328226
rect 387594 328170 387662 328226
rect 387718 328170 387786 328226
rect 387842 328170 387866 328226
rect 387390 328102 387866 328170
rect 387390 328046 387414 328102
rect 387470 328046 387538 328102
rect 387594 328046 387662 328102
rect 387718 328046 387786 328102
rect 387842 328046 387866 328102
rect 387390 327978 387866 328046
rect 387390 327922 387414 327978
rect 387470 327922 387538 327978
rect 387594 327922 387662 327978
rect 387718 327922 387786 327978
rect 387842 327922 387866 327978
rect 387390 327888 387866 327922
rect 377778 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 378398 316350
rect 377778 316226 378398 316294
rect 377778 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 378398 316226
rect 377778 316102 378398 316170
rect 377778 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 378398 316102
rect 377778 315978 378398 316046
rect 377778 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 378398 315978
rect 377778 298350 378398 315922
rect 386590 316350 387066 316384
rect 386590 316294 386614 316350
rect 386670 316294 386738 316350
rect 386794 316294 386862 316350
rect 386918 316294 386986 316350
rect 387042 316294 387066 316350
rect 386590 316226 387066 316294
rect 386590 316170 386614 316226
rect 386670 316170 386738 316226
rect 386794 316170 386862 316226
rect 386918 316170 386986 316226
rect 387042 316170 387066 316226
rect 386590 316102 387066 316170
rect 386590 316046 386614 316102
rect 386670 316046 386738 316102
rect 386794 316046 386862 316102
rect 386918 316046 386986 316102
rect 387042 316046 387066 316102
rect 386590 315978 387066 316046
rect 386590 315922 386614 315978
rect 386670 315922 386738 315978
rect 386794 315922 386862 315978
rect 386918 315922 386986 315978
rect 387042 315922 387066 315978
rect 386590 315888 387066 315922
rect 387390 310350 387866 310384
rect 387390 310294 387414 310350
rect 387470 310294 387538 310350
rect 387594 310294 387662 310350
rect 387718 310294 387786 310350
rect 387842 310294 387866 310350
rect 387390 310226 387866 310294
rect 387390 310170 387414 310226
rect 387470 310170 387538 310226
rect 387594 310170 387662 310226
rect 387718 310170 387786 310226
rect 387842 310170 387866 310226
rect 387390 310102 387866 310170
rect 387390 310046 387414 310102
rect 387470 310046 387538 310102
rect 387594 310046 387662 310102
rect 387718 310046 387786 310102
rect 387842 310046 387866 310102
rect 387390 309978 387866 310046
rect 387390 309922 387414 309978
rect 387470 309922 387538 309978
rect 387594 309922 387662 309978
rect 387718 309922 387786 309978
rect 387842 309922 387866 309978
rect 387390 309888 387866 309922
rect 388108 302372 388164 302382
rect 387996 302316 388108 302338
rect 387996 302282 388164 302316
rect 387996 301798 388052 302282
rect 387996 301732 388052 301742
rect 387996 300692 388164 300718
rect 387996 300662 388108 300692
rect 387996 300358 388052 300662
rect 388108 300626 388164 300636
rect 387996 300292 388052 300302
rect 388220 300580 388276 300590
rect 388220 300358 388276 300524
rect 388220 300292 388276 300302
rect 377778 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 378398 298350
rect 377778 298226 378398 298294
rect 377778 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 378398 298226
rect 377778 298102 378398 298170
rect 377778 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 378398 298102
rect 377778 297978 378398 298046
rect 377778 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 378398 297978
rect 377778 280350 378398 297922
rect 386590 298350 387066 298384
rect 386590 298294 386614 298350
rect 386670 298294 386738 298350
rect 386794 298294 386862 298350
rect 386918 298294 386986 298350
rect 387042 298294 387066 298350
rect 386590 298226 387066 298294
rect 386590 298170 386614 298226
rect 386670 298170 386738 298226
rect 386794 298170 386862 298226
rect 386918 298170 386986 298226
rect 387042 298170 387066 298226
rect 386590 298102 387066 298170
rect 386590 298046 386614 298102
rect 386670 298046 386738 298102
rect 386794 298046 386862 298102
rect 386918 298046 386986 298102
rect 387042 298046 387066 298102
rect 386590 297978 387066 298046
rect 386590 297922 386614 297978
rect 386670 297922 386738 297978
rect 386794 297922 386862 297978
rect 386918 297922 386986 297978
rect 387042 297922 387066 297978
rect 386590 297888 387066 297922
rect 388220 297332 388276 297342
rect 388220 296938 388276 297276
rect 387996 296882 388276 296938
rect 388444 297220 388500 297230
rect 388444 296938 388500 297164
rect 390572 297118 390628 328524
rect 390572 297052 390628 297062
rect 404778 328350 405398 345922
rect 404778 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 405398 328350
rect 404778 328226 405398 328294
rect 404778 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 405398 328226
rect 404778 328102 405398 328170
rect 404778 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 405398 328102
rect 404778 327978 405398 328046
rect 404778 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 405398 327978
rect 404778 310350 405398 327922
rect 404778 310294 404874 310350
rect 404930 310294 404998 310350
rect 405054 310294 405122 310350
rect 405178 310294 405246 310350
rect 405302 310294 405398 310350
rect 404778 310226 405398 310294
rect 404778 310170 404874 310226
rect 404930 310170 404998 310226
rect 405054 310170 405122 310226
rect 405178 310170 405246 310226
rect 405302 310170 405398 310226
rect 404778 310102 405398 310170
rect 404778 310046 404874 310102
rect 404930 310046 404998 310102
rect 405054 310046 405122 310102
rect 405178 310046 405246 310102
rect 405302 310046 405398 310102
rect 404778 309978 405398 310046
rect 404778 309922 404874 309978
rect 404930 309922 404998 309978
rect 405054 309922 405122 309978
rect 405178 309922 405246 309978
rect 405302 309922 405398 309978
rect 387996 296758 388052 296882
rect 388444 296872 388500 296882
rect 387996 296692 388052 296702
rect 387390 292350 387866 292384
rect 387390 292294 387414 292350
rect 387470 292294 387538 292350
rect 387594 292294 387662 292350
rect 387718 292294 387786 292350
rect 387842 292294 387866 292350
rect 404778 292350 405398 309922
rect 387390 292226 387866 292294
rect 388108 292292 388164 292302
rect 387390 292170 387414 292226
rect 387470 292170 387538 292226
rect 387594 292170 387662 292226
rect 387718 292170 387786 292226
rect 387842 292170 387866 292226
rect 387390 292102 387866 292170
rect 387390 292046 387414 292102
rect 387470 292046 387538 292102
rect 387594 292046 387662 292102
rect 387718 292046 387786 292102
rect 387842 292046 387866 292102
rect 387390 291978 387866 292046
rect 387390 291922 387414 291978
rect 387470 291922 387538 291978
rect 387594 291922 387662 291978
rect 387718 291922 387786 291978
rect 387842 291922 387866 291978
rect 387390 291888 387866 291922
rect 387996 292236 388108 292258
rect 387996 292202 388164 292236
rect 404778 292294 404874 292350
rect 404930 292294 404998 292350
rect 405054 292294 405122 292350
rect 405178 292294 405246 292350
rect 405302 292294 405398 292350
rect 404778 292226 405398 292294
rect 387996 291718 388052 292202
rect 387996 291652 388052 291662
rect 404778 292170 404874 292226
rect 404930 292170 404998 292226
rect 405054 292170 405122 292226
rect 405178 292170 405246 292226
rect 405302 292170 405398 292226
rect 404778 292102 405398 292170
rect 404778 292046 404874 292102
rect 404930 292046 404998 292102
rect 405054 292046 405122 292102
rect 405178 292046 405246 292102
rect 405302 292046 405398 292102
rect 404778 291978 405398 292046
rect 404778 291922 404874 291978
rect 404930 291922 404998 291978
rect 405054 291922 405122 291978
rect 405178 291922 405246 291978
rect 405302 291922 405398 291978
rect 387996 290612 388164 290638
rect 387996 290582 388108 290612
rect 387996 290278 388052 290582
rect 388108 290546 388164 290556
rect 387996 290212 388052 290222
rect 377778 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 378398 280350
rect 377778 280226 378398 280294
rect 377778 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 378398 280226
rect 377778 280102 378398 280170
rect 377778 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 378398 280102
rect 377778 279978 378398 280046
rect 377778 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 378398 279978
rect 377778 262350 378398 279922
rect 377778 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 378398 262350
rect 377778 262226 378398 262294
rect 377778 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 378398 262226
rect 377778 262102 378398 262170
rect 377778 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 378398 262102
rect 377778 261978 378398 262046
rect 377778 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 378398 261978
rect 375004 259140 375060 259150
rect 374058 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 374678 256350
rect 374058 256226 374678 256294
rect 374058 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 374678 256226
rect 374058 256102 374678 256170
rect 374058 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 374678 256102
rect 374058 255978 374678 256046
rect 374058 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 374678 255978
rect 374058 238350 374678 255922
rect 374892 258692 374948 258702
rect 374892 243628 374948 258636
rect 375004 255388 375060 259084
rect 375004 255332 375172 255388
rect 374058 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 374678 238350
rect 374058 238226 374678 238294
rect 374058 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 374678 238226
rect 374058 238102 374678 238170
rect 374058 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 374678 238102
rect 374058 237978 374678 238046
rect 374058 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 374678 237978
rect 374058 220350 374678 237922
rect 374058 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 374678 220350
rect 374058 220226 374678 220294
rect 374058 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 374678 220226
rect 374058 220102 374678 220170
rect 374058 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 374678 220102
rect 374058 219978 374678 220046
rect 374058 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 374678 219978
rect 374058 202350 374678 219922
rect 374058 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 374678 202350
rect 374058 202226 374678 202294
rect 374058 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 374678 202226
rect 374058 202102 374678 202170
rect 374058 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 374678 202102
rect 374058 201978 374678 202046
rect 374058 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 374678 201978
rect 374058 184350 374678 201922
rect 374058 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 374678 184350
rect 374058 184226 374678 184294
rect 374058 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 374678 184226
rect 374058 184102 374678 184170
rect 374058 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 374678 184102
rect 374058 183978 374678 184046
rect 374058 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 374678 183978
rect 374058 166350 374678 183922
rect 374058 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 374678 166350
rect 374058 166226 374678 166294
rect 374058 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 374678 166226
rect 374058 166102 374678 166170
rect 374058 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 374678 166102
rect 374058 165978 374678 166046
rect 374058 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 374678 165978
rect 374058 148350 374678 165922
rect 374058 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 374678 148350
rect 374058 148226 374678 148294
rect 374058 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 374678 148226
rect 374058 148102 374678 148170
rect 374058 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 374678 148102
rect 374058 147978 374678 148046
rect 374058 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 374678 147978
rect 361106 130350 361582 130384
rect 361106 130294 361130 130350
rect 361186 130294 361254 130350
rect 361310 130294 361378 130350
rect 361434 130294 361502 130350
rect 361558 130294 361582 130350
rect 361106 130226 361582 130294
rect 361106 130170 361130 130226
rect 361186 130170 361254 130226
rect 361310 130170 361378 130226
rect 361434 130170 361502 130226
rect 361558 130170 361582 130226
rect 361106 130102 361582 130170
rect 361106 130046 361130 130102
rect 361186 130046 361254 130102
rect 361310 130046 361378 130102
rect 361434 130046 361502 130102
rect 361558 130046 361582 130102
rect 361106 129978 361582 130046
rect 361106 129922 361130 129978
rect 361186 129922 361254 129978
rect 361310 129922 361378 129978
rect 361434 129922 361502 129978
rect 361558 129922 361582 129978
rect 361106 129888 361582 129922
rect 374058 130350 374678 147922
rect 374780 243572 374948 243628
rect 374780 141428 374836 243572
rect 375116 142548 375172 255332
rect 375116 141876 375172 142492
rect 375116 141810 375172 141820
rect 377778 244350 378398 261922
rect 404778 274350 405398 291922
rect 404778 274294 404874 274350
rect 404930 274294 404998 274350
rect 405054 274294 405122 274350
rect 405178 274294 405246 274350
rect 405302 274294 405398 274350
rect 404778 274226 405398 274294
rect 404778 274170 404874 274226
rect 404930 274170 404998 274226
rect 405054 274170 405122 274226
rect 405178 274170 405246 274226
rect 405302 274170 405398 274226
rect 404778 274102 405398 274170
rect 404778 274046 404874 274102
rect 404930 274046 404998 274102
rect 405054 274046 405122 274102
rect 405178 274046 405246 274102
rect 405302 274046 405398 274102
rect 404778 273978 405398 274046
rect 404778 273922 404874 273978
rect 404930 273922 404998 273978
rect 405054 273922 405122 273978
rect 405178 273922 405246 273978
rect 405302 273922 405398 273978
rect 385756 259140 385812 259150
rect 385420 258916 385476 258926
rect 385420 255388 385476 258860
rect 385420 255332 385588 255388
rect 377778 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 378398 244350
rect 377778 244226 378398 244294
rect 377778 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 378398 244226
rect 377778 244102 378398 244170
rect 377778 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 378398 244102
rect 377778 243978 378398 244046
rect 377778 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 378398 243978
rect 377778 226350 378398 243922
rect 377778 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 378398 226350
rect 377778 226226 378398 226294
rect 377778 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 378398 226226
rect 377778 226102 378398 226170
rect 377778 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 378398 226102
rect 377778 225978 378398 226046
rect 377778 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 378398 225978
rect 377778 208350 378398 225922
rect 377778 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208294 378398 208350
rect 377778 208226 378398 208294
rect 377778 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208170 378398 208226
rect 377778 208102 378398 208170
rect 377778 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 378398 208102
rect 377778 207978 378398 208046
rect 377778 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 378398 207978
rect 377778 190350 378398 207922
rect 377778 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 378398 190350
rect 377778 190226 378398 190294
rect 377778 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 378398 190226
rect 377778 190102 378398 190170
rect 377778 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 378398 190102
rect 377778 189978 378398 190046
rect 377778 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 378398 189978
rect 377778 172350 378398 189922
rect 377778 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 378398 172350
rect 377778 172226 378398 172294
rect 377778 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 378398 172226
rect 377778 172102 378398 172170
rect 377778 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 378398 172102
rect 377778 171978 378398 172046
rect 377778 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 378398 171978
rect 377778 154350 378398 171922
rect 377778 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 378398 154350
rect 377778 154226 378398 154294
rect 377778 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 378398 154226
rect 377778 154102 378398 154170
rect 377778 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 378398 154102
rect 377778 153978 378398 154046
rect 377778 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 378398 153978
rect 374780 141362 374836 141372
rect 374058 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 374678 130350
rect 374058 130226 374678 130294
rect 374058 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 374678 130226
rect 374058 130102 374678 130170
rect 374058 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 374678 130102
rect 374058 129978 374678 130046
rect 374058 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 374678 129978
rect 361906 118350 362382 118384
rect 361906 118294 361930 118350
rect 361986 118294 362054 118350
rect 362110 118294 362178 118350
rect 362234 118294 362302 118350
rect 362358 118294 362382 118350
rect 361906 118226 362382 118294
rect 361906 118170 361930 118226
rect 361986 118170 362054 118226
rect 362110 118170 362178 118226
rect 362234 118170 362302 118226
rect 362358 118170 362382 118226
rect 361906 118102 362382 118170
rect 361906 118046 361930 118102
rect 361986 118046 362054 118102
rect 362110 118046 362178 118102
rect 362234 118046 362302 118102
rect 362358 118046 362382 118102
rect 361906 117978 362382 118046
rect 361906 117922 361930 117978
rect 361986 117922 362054 117978
rect 362110 117922 362178 117978
rect 362234 117922 362302 117978
rect 362358 117922 362382 117978
rect 361906 117888 362382 117922
rect 361106 112350 361582 112384
rect 361106 112294 361130 112350
rect 361186 112294 361254 112350
rect 361310 112294 361378 112350
rect 361434 112294 361502 112350
rect 361558 112294 361582 112350
rect 361106 112226 361582 112294
rect 361106 112170 361130 112226
rect 361186 112170 361254 112226
rect 361310 112170 361378 112226
rect 361434 112170 361502 112226
rect 361558 112170 361582 112226
rect 361106 112102 361582 112170
rect 361106 112046 361130 112102
rect 361186 112046 361254 112102
rect 361310 112046 361378 112102
rect 361434 112046 361502 112102
rect 361558 112046 361582 112102
rect 361106 111978 361582 112046
rect 361106 111922 361130 111978
rect 361186 111922 361254 111978
rect 361310 111922 361378 111978
rect 361434 111922 361502 111978
rect 361558 111922 361582 111978
rect 361106 111888 361582 111922
rect 374058 112350 374678 129922
rect 374058 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 374678 112350
rect 374058 112226 374678 112294
rect 374058 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 374678 112226
rect 374058 112102 374678 112170
rect 374058 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 374678 112102
rect 374058 111978 374678 112046
rect 374058 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 374678 111978
rect 361906 100350 362382 100384
rect 361906 100294 361930 100350
rect 361986 100294 362054 100350
rect 362110 100294 362178 100350
rect 362234 100294 362302 100350
rect 362358 100294 362382 100350
rect 361906 100226 362382 100294
rect 361906 100170 361930 100226
rect 361986 100170 362054 100226
rect 362110 100170 362178 100226
rect 362234 100170 362302 100226
rect 362358 100170 362382 100226
rect 361906 100102 362382 100170
rect 361906 100046 361930 100102
rect 361986 100046 362054 100102
rect 362110 100046 362178 100102
rect 362234 100046 362302 100102
rect 362358 100046 362382 100102
rect 361906 99978 362382 100046
rect 361906 99922 361930 99978
rect 361986 99922 362054 99978
rect 362110 99922 362178 99978
rect 362234 99922 362302 99978
rect 362358 99922 362382 99978
rect 361906 99888 362382 99922
rect 361106 94350 361582 94384
rect 361106 94294 361130 94350
rect 361186 94294 361254 94350
rect 361310 94294 361378 94350
rect 361434 94294 361502 94350
rect 361558 94294 361582 94350
rect 361106 94226 361582 94294
rect 361106 94170 361130 94226
rect 361186 94170 361254 94226
rect 361310 94170 361378 94226
rect 361434 94170 361502 94226
rect 361558 94170 361582 94226
rect 361106 94102 361582 94170
rect 361106 94046 361130 94102
rect 361186 94046 361254 94102
rect 361310 94046 361378 94102
rect 361434 94046 361502 94102
rect 361558 94046 361582 94102
rect 361106 93978 361582 94046
rect 361106 93922 361130 93978
rect 361186 93922 361254 93978
rect 361310 93922 361378 93978
rect 361434 93922 361502 93978
rect 361558 93922 361582 93978
rect 361106 93888 361582 93922
rect 374058 94350 374678 111922
rect 374058 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 374678 94350
rect 374058 94226 374678 94294
rect 374058 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 374678 94226
rect 374058 94102 374678 94170
rect 374058 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 374678 94102
rect 374058 93978 374678 94046
rect 374058 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 374678 93978
rect 361906 82350 362382 82384
rect 361906 82294 361930 82350
rect 361986 82294 362054 82350
rect 362110 82294 362178 82350
rect 362234 82294 362302 82350
rect 362358 82294 362382 82350
rect 361906 82226 362382 82294
rect 361906 82170 361930 82226
rect 361986 82170 362054 82226
rect 362110 82170 362178 82226
rect 362234 82170 362302 82226
rect 362358 82170 362382 82226
rect 361906 82102 362382 82170
rect 361906 82046 361930 82102
rect 361986 82046 362054 82102
rect 362110 82046 362178 82102
rect 362234 82046 362302 82102
rect 362358 82046 362382 82102
rect 361906 81978 362382 82046
rect 361906 81922 361930 81978
rect 361986 81922 362054 81978
rect 362110 81922 362178 81978
rect 362234 81922 362302 81978
rect 362358 81922 362382 81978
rect 361906 81888 362382 81922
rect 361106 76350 361582 76384
rect 361106 76294 361130 76350
rect 361186 76294 361254 76350
rect 361310 76294 361378 76350
rect 361434 76294 361502 76350
rect 361558 76294 361582 76350
rect 361106 76226 361582 76294
rect 361106 76170 361130 76226
rect 361186 76170 361254 76226
rect 361310 76170 361378 76226
rect 361434 76170 361502 76226
rect 361558 76170 361582 76226
rect 361106 76102 361582 76170
rect 361106 76046 361130 76102
rect 361186 76046 361254 76102
rect 361310 76046 361378 76102
rect 361434 76046 361502 76102
rect 361558 76046 361582 76102
rect 361106 75978 361582 76046
rect 361106 75922 361130 75978
rect 361186 75922 361254 75978
rect 361310 75922 361378 75978
rect 361434 75922 361502 75978
rect 361558 75922 361582 75978
rect 361106 75888 361582 75922
rect 374058 76350 374678 93922
rect 374058 76294 374154 76350
rect 374210 76294 374278 76350
rect 374334 76294 374402 76350
rect 374458 76294 374526 76350
rect 374582 76294 374678 76350
rect 374058 76226 374678 76294
rect 374058 76170 374154 76226
rect 374210 76170 374278 76226
rect 374334 76170 374402 76226
rect 374458 76170 374526 76226
rect 374582 76170 374678 76226
rect 374058 76102 374678 76170
rect 374058 76046 374154 76102
rect 374210 76046 374278 76102
rect 374334 76046 374402 76102
rect 374458 76046 374526 76102
rect 374582 76046 374678 76102
rect 374058 75978 374678 76046
rect 374058 75922 374154 75978
rect 374210 75922 374278 75978
rect 374334 75922 374402 75978
rect 374458 75922 374526 75978
rect 374582 75922 374678 75978
rect 361906 64350 362382 64384
rect 361906 64294 361930 64350
rect 361986 64294 362054 64350
rect 362110 64294 362178 64350
rect 362234 64294 362302 64350
rect 362358 64294 362382 64350
rect 361906 64226 362382 64294
rect 361906 64170 361930 64226
rect 361986 64170 362054 64226
rect 362110 64170 362178 64226
rect 362234 64170 362302 64226
rect 362358 64170 362382 64226
rect 361906 64102 362382 64170
rect 361906 64046 361930 64102
rect 361986 64046 362054 64102
rect 362110 64046 362178 64102
rect 362234 64046 362302 64102
rect 362358 64046 362382 64102
rect 361906 63978 362382 64046
rect 361906 63922 361930 63978
rect 361986 63922 362054 63978
rect 362110 63922 362178 63978
rect 362234 63922 362302 63978
rect 362358 63922 362382 63978
rect 361906 63888 362382 63922
rect 361106 58350 361582 58384
rect 361106 58294 361130 58350
rect 361186 58294 361254 58350
rect 361310 58294 361378 58350
rect 361434 58294 361502 58350
rect 361558 58294 361582 58350
rect 361106 58226 361582 58294
rect 361106 58170 361130 58226
rect 361186 58170 361254 58226
rect 361310 58170 361378 58226
rect 361434 58170 361502 58226
rect 361558 58170 361582 58226
rect 361106 58102 361582 58170
rect 361106 58046 361130 58102
rect 361186 58046 361254 58102
rect 361310 58046 361378 58102
rect 361434 58046 361502 58102
rect 361558 58046 361582 58102
rect 361106 57978 361582 58046
rect 361106 57922 361130 57978
rect 361186 57922 361254 57978
rect 361310 57922 361378 57978
rect 361434 57922 361502 57978
rect 361558 57922 361582 57978
rect 361106 57888 361582 57922
rect 374058 58350 374678 75922
rect 374058 58294 374154 58350
rect 374210 58294 374278 58350
rect 374334 58294 374402 58350
rect 374458 58294 374526 58350
rect 374582 58294 374678 58350
rect 374058 58226 374678 58294
rect 374058 58170 374154 58226
rect 374210 58170 374278 58226
rect 374334 58170 374402 58226
rect 374458 58170 374526 58226
rect 374582 58170 374678 58226
rect 374058 58102 374678 58170
rect 374058 58046 374154 58102
rect 374210 58046 374278 58102
rect 374334 58046 374402 58102
rect 374458 58046 374526 58102
rect 374582 58046 374678 58102
rect 374058 57978 374678 58046
rect 374058 57922 374154 57978
rect 374210 57922 374278 57978
rect 374334 57922 374402 57978
rect 374458 57922 374526 57978
rect 374582 57922 374678 57978
rect 361906 46350 362382 46384
rect 361906 46294 361930 46350
rect 361986 46294 362054 46350
rect 362110 46294 362178 46350
rect 362234 46294 362302 46350
rect 362358 46294 362382 46350
rect 361906 46226 362382 46294
rect 361906 46170 361930 46226
rect 361986 46170 362054 46226
rect 362110 46170 362178 46226
rect 362234 46170 362302 46226
rect 362358 46170 362382 46226
rect 361906 46102 362382 46170
rect 361906 46046 361930 46102
rect 361986 46046 362054 46102
rect 362110 46046 362178 46102
rect 362234 46046 362302 46102
rect 362358 46046 362382 46102
rect 361906 45978 362382 46046
rect 361906 45922 361930 45978
rect 361986 45922 362054 45978
rect 362110 45922 362178 45978
rect 362234 45922 362302 45978
rect 362358 45922 362382 45978
rect 361906 45888 362382 45922
rect 360332 4498 360388 4508
rect 374058 40350 374678 57922
rect 374058 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 374678 40350
rect 374058 40226 374678 40294
rect 374058 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 374678 40226
rect 374058 40102 374678 40170
rect 374058 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 374678 40102
rect 374058 39978 374678 40046
rect 374058 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 374678 39978
rect 374058 22350 374678 39922
rect 374058 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 374678 22350
rect 374058 22226 374678 22294
rect 374058 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 374678 22226
rect 374058 22102 374678 22170
rect 374058 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 374678 22102
rect 374058 21978 374678 22046
rect 374058 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 374678 21978
rect 358652 4162 358708 4172
rect 374058 4350 374678 21922
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 347058 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 347678 -1120
rect 347058 -1244 347678 -1176
rect 347058 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 347678 -1244
rect 347058 -1368 347678 -1300
rect 347058 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 347678 -1368
rect 347058 -1492 347678 -1424
rect 347058 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 347678 -1492
rect 347058 -1644 347678 -1548
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 377778 136350 378398 153922
rect 385532 142660 385588 255332
rect 385532 141316 385588 142604
rect 385532 141250 385588 141260
rect 385756 140420 385812 259084
rect 385756 139860 385812 140364
rect 390572 259140 390628 259150
rect 390572 139972 390628 259084
rect 393932 259140 393988 259150
rect 392252 259028 392308 259038
rect 392252 140868 392308 258972
rect 392252 140802 392308 140812
rect 392476 259028 392532 259038
rect 392476 140532 392532 258972
rect 393932 140756 393988 259084
rect 393932 140690 393988 140700
rect 397292 259140 397348 259150
rect 392476 140466 392532 140476
rect 390572 139906 390628 139916
rect 385756 139794 385812 139804
rect 397292 138852 397348 259084
rect 397292 138786 397348 138796
rect 404778 256350 405398 273922
rect 404778 256294 404874 256350
rect 404930 256294 404998 256350
rect 405054 256294 405122 256350
rect 405178 256294 405246 256350
rect 405302 256294 405398 256350
rect 404778 256226 405398 256294
rect 404778 256170 404874 256226
rect 404930 256170 404998 256226
rect 405054 256170 405122 256226
rect 405178 256170 405246 256226
rect 405302 256170 405398 256226
rect 404778 256102 405398 256170
rect 404778 256046 404874 256102
rect 404930 256046 404998 256102
rect 405054 256046 405122 256102
rect 405178 256046 405246 256102
rect 405302 256046 405398 256102
rect 404778 255978 405398 256046
rect 404778 255922 404874 255978
rect 404930 255922 404998 255978
rect 405054 255922 405122 255978
rect 405178 255922 405246 255978
rect 405302 255922 405398 255978
rect 404778 238350 405398 255922
rect 404778 238294 404874 238350
rect 404930 238294 404998 238350
rect 405054 238294 405122 238350
rect 405178 238294 405246 238350
rect 405302 238294 405398 238350
rect 404778 238226 405398 238294
rect 404778 238170 404874 238226
rect 404930 238170 404998 238226
rect 405054 238170 405122 238226
rect 405178 238170 405246 238226
rect 405302 238170 405398 238226
rect 404778 238102 405398 238170
rect 404778 238046 404874 238102
rect 404930 238046 404998 238102
rect 405054 238046 405122 238102
rect 405178 238046 405246 238102
rect 405302 238046 405398 238102
rect 404778 237978 405398 238046
rect 404778 237922 404874 237978
rect 404930 237922 404998 237978
rect 405054 237922 405122 237978
rect 405178 237922 405246 237978
rect 405302 237922 405398 237978
rect 404778 220350 405398 237922
rect 404778 220294 404874 220350
rect 404930 220294 404998 220350
rect 405054 220294 405122 220350
rect 405178 220294 405246 220350
rect 405302 220294 405398 220350
rect 404778 220226 405398 220294
rect 404778 220170 404874 220226
rect 404930 220170 404998 220226
rect 405054 220170 405122 220226
rect 405178 220170 405246 220226
rect 405302 220170 405398 220226
rect 404778 220102 405398 220170
rect 404778 220046 404874 220102
rect 404930 220046 404998 220102
rect 405054 220046 405122 220102
rect 405178 220046 405246 220102
rect 405302 220046 405398 220102
rect 404778 219978 405398 220046
rect 404778 219922 404874 219978
rect 404930 219922 404998 219978
rect 405054 219922 405122 219978
rect 405178 219922 405246 219978
rect 405302 219922 405398 219978
rect 404778 202350 405398 219922
rect 404778 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 405398 202350
rect 404778 202226 405398 202294
rect 404778 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 405398 202226
rect 404778 202102 405398 202170
rect 404778 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 405398 202102
rect 404778 201978 405398 202046
rect 404778 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 405398 201978
rect 404778 184350 405398 201922
rect 404778 184294 404874 184350
rect 404930 184294 404998 184350
rect 405054 184294 405122 184350
rect 405178 184294 405246 184350
rect 405302 184294 405398 184350
rect 404778 184226 405398 184294
rect 404778 184170 404874 184226
rect 404930 184170 404998 184226
rect 405054 184170 405122 184226
rect 405178 184170 405246 184226
rect 405302 184170 405398 184226
rect 404778 184102 405398 184170
rect 404778 184046 404874 184102
rect 404930 184046 404998 184102
rect 405054 184046 405122 184102
rect 405178 184046 405246 184102
rect 405302 184046 405398 184102
rect 404778 183978 405398 184046
rect 404778 183922 404874 183978
rect 404930 183922 404998 183978
rect 405054 183922 405122 183978
rect 405178 183922 405246 183978
rect 405302 183922 405398 183978
rect 404778 166350 405398 183922
rect 404778 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 405398 166350
rect 404778 166226 405398 166294
rect 404778 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 405398 166226
rect 404778 166102 405398 166170
rect 404778 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 405398 166102
rect 404778 165978 405398 166046
rect 404778 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 405398 165978
rect 404778 148350 405398 165922
rect 404778 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 405398 148350
rect 404778 148226 405398 148294
rect 404778 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 405398 148226
rect 404778 148102 405398 148170
rect 404778 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 405398 148102
rect 404778 147978 405398 148046
rect 404778 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 405398 147978
rect 377778 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 378398 136350
rect 377778 136226 378398 136294
rect 377778 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 378398 136226
rect 377778 136102 378398 136170
rect 377778 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 378398 136102
rect 377778 135978 378398 136046
rect 377778 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 378398 135978
rect 377778 118350 378398 135922
rect 377778 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 378398 118350
rect 377778 118226 378398 118294
rect 377778 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 378398 118226
rect 377778 118102 378398 118170
rect 377778 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 378398 118102
rect 377778 117978 378398 118046
rect 377778 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 378398 117978
rect 377778 100350 378398 117922
rect 377778 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 378398 100350
rect 377778 100226 378398 100294
rect 377778 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 378398 100226
rect 377778 100102 378398 100170
rect 377778 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 378398 100102
rect 377778 99978 378398 100046
rect 377778 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 378398 99978
rect 377778 82350 378398 99922
rect 377778 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 378398 82350
rect 377778 82226 378398 82294
rect 377778 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 378398 82226
rect 377778 82102 378398 82170
rect 377778 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 378398 82102
rect 377778 81978 378398 82046
rect 377778 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 378398 81978
rect 377778 64350 378398 81922
rect 377778 64294 377874 64350
rect 377930 64294 377998 64350
rect 378054 64294 378122 64350
rect 378178 64294 378246 64350
rect 378302 64294 378398 64350
rect 377778 64226 378398 64294
rect 377778 64170 377874 64226
rect 377930 64170 377998 64226
rect 378054 64170 378122 64226
rect 378178 64170 378246 64226
rect 378302 64170 378398 64226
rect 377778 64102 378398 64170
rect 377778 64046 377874 64102
rect 377930 64046 377998 64102
rect 378054 64046 378122 64102
rect 378178 64046 378246 64102
rect 378302 64046 378398 64102
rect 377778 63978 378398 64046
rect 377778 63922 377874 63978
rect 377930 63922 377998 63978
rect 378054 63922 378122 63978
rect 378178 63922 378246 63978
rect 378302 63922 378398 63978
rect 377778 46350 378398 63922
rect 377778 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 378398 46350
rect 377778 46226 378398 46294
rect 377778 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 378398 46226
rect 377778 46102 378398 46170
rect 377778 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 378398 46102
rect 377778 45978 378398 46046
rect 377778 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 378398 45978
rect 377778 28350 378398 45922
rect 377778 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 378398 28350
rect 377778 28226 378398 28294
rect 377778 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 378398 28226
rect 377778 28102 378398 28170
rect 377778 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 378398 28102
rect 377778 27978 378398 28046
rect 377778 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 378398 27978
rect 377778 10350 378398 27922
rect 377778 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 378398 10350
rect 377778 10226 378398 10294
rect 377778 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 378398 10226
rect 377778 10102 378398 10170
rect 377778 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 378398 10102
rect 377778 9978 378398 10046
rect 377778 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 378398 9978
rect 377778 -1120 378398 9922
rect 377778 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 378398 -1120
rect 377778 -1244 378398 -1176
rect 377778 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 378398 -1244
rect 377778 -1368 378398 -1300
rect 377778 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 378398 -1368
rect 377778 -1492 378398 -1424
rect 377778 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 378398 -1492
rect 377778 -1644 378398 -1548
rect 404778 130350 405398 147922
rect 404778 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 405398 130350
rect 404778 130226 405398 130294
rect 404778 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 405398 130226
rect 404778 130102 405398 130170
rect 404778 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 405398 130102
rect 404778 129978 405398 130046
rect 404778 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 405398 129978
rect 404778 112350 405398 129922
rect 404778 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 405398 112350
rect 404778 112226 405398 112294
rect 404778 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 405398 112226
rect 404778 112102 405398 112170
rect 404778 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 405398 112102
rect 404778 111978 405398 112046
rect 404778 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 405398 111978
rect 404778 94350 405398 111922
rect 404778 94294 404874 94350
rect 404930 94294 404998 94350
rect 405054 94294 405122 94350
rect 405178 94294 405246 94350
rect 405302 94294 405398 94350
rect 404778 94226 405398 94294
rect 404778 94170 404874 94226
rect 404930 94170 404998 94226
rect 405054 94170 405122 94226
rect 405178 94170 405246 94226
rect 405302 94170 405398 94226
rect 404778 94102 405398 94170
rect 404778 94046 404874 94102
rect 404930 94046 404998 94102
rect 405054 94046 405122 94102
rect 405178 94046 405246 94102
rect 405302 94046 405398 94102
rect 404778 93978 405398 94046
rect 404778 93922 404874 93978
rect 404930 93922 404998 93978
rect 405054 93922 405122 93978
rect 405178 93922 405246 93978
rect 405302 93922 405398 93978
rect 404778 76350 405398 93922
rect 404778 76294 404874 76350
rect 404930 76294 404998 76350
rect 405054 76294 405122 76350
rect 405178 76294 405246 76350
rect 405302 76294 405398 76350
rect 404778 76226 405398 76294
rect 404778 76170 404874 76226
rect 404930 76170 404998 76226
rect 405054 76170 405122 76226
rect 405178 76170 405246 76226
rect 405302 76170 405398 76226
rect 404778 76102 405398 76170
rect 404778 76046 404874 76102
rect 404930 76046 404998 76102
rect 405054 76046 405122 76102
rect 405178 76046 405246 76102
rect 405302 76046 405398 76102
rect 404778 75978 405398 76046
rect 404778 75922 404874 75978
rect 404930 75922 404998 75978
rect 405054 75922 405122 75978
rect 405178 75922 405246 75978
rect 405302 75922 405398 75978
rect 404778 58350 405398 75922
rect 404778 58294 404874 58350
rect 404930 58294 404998 58350
rect 405054 58294 405122 58350
rect 405178 58294 405246 58350
rect 405302 58294 405398 58350
rect 404778 58226 405398 58294
rect 404778 58170 404874 58226
rect 404930 58170 404998 58226
rect 405054 58170 405122 58226
rect 405178 58170 405246 58226
rect 405302 58170 405398 58226
rect 404778 58102 405398 58170
rect 404778 58046 404874 58102
rect 404930 58046 404998 58102
rect 405054 58046 405122 58102
rect 405178 58046 405246 58102
rect 405302 58046 405398 58102
rect 404778 57978 405398 58046
rect 404778 57922 404874 57978
rect 404930 57922 404998 57978
rect 405054 57922 405122 57978
rect 405178 57922 405246 57978
rect 405302 57922 405398 57978
rect 404778 40350 405398 57922
rect 404778 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 405398 40350
rect 404778 40226 405398 40294
rect 404778 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 405398 40226
rect 404778 40102 405398 40170
rect 404778 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 405398 40102
rect 404778 39978 405398 40046
rect 404778 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 405398 39978
rect 404778 22350 405398 39922
rect 404778 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 405398 22350
rect 404778 22226 405398 22294
rect 404778 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 405398 22226
rect 404778 22102 405398 22170
rect 404778 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 405398 22102
rect 404778 21978 405398 22046
rect 404778 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 405398 21978
rect 404778 4350 405398 21922
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 408498 388350 409118 402722
rect 408498 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388294 409118 388350
rect 408498 388226 409118 388294
rect 408498 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 409118 388226
rect 408498 388102 409118 388170
rect 408498 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 409118 388102
rect 408498 387978 409118 388046
rect 408498 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 409118 387978
rect 408498 370350 409118 387922
rect 408498 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 409118 370350
rect 408498 370226 409118 370294
rect 408498 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 409118 370226
rect 408498 370102 409118 370170
rect 408498 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 409118 370102
rect 408498 369978 409118 370046
rect 408498 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 409118 369978
rect 408498 352350 409118 369922
rect 408498 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 409118 352350
rect 408498 352226 409118 352294
rect 408498 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 409118 352226
rect 408498 352102 409118 352170
rect 408498 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 409118 352102
rect 408498 351978 409118 352046
rect 408498 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 409118 351978
rect 408498 334350 409118 351922
rect 408498 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 409118 334350
rect 408498 334226 409118 334294
rect 408498 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 409118 334226
rect 408498 334102 409118 334170
rect 408498 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 409118 334102
rect 408498 333978 409118 334046
rect 408498 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 409118 333978
rect 408498 316350 409118 333922
rect 408498 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 409118 316350
rect 408498 316226 409118 316294
rect 408498 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 409118 316226
rect 408498 316102 409118 316170
rect 408498 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 409118 316102
rect 408498 315978 409118 316046
rect 408498 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 409118 315978
rect 408498 298350 409118 315922
rect 408498 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 409118 298350
rect 408498 298226 409118 298294
rect 408498 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 409118 298226
rect 408498 298102 409118 298170
rect 408498 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 409118 298102
rect 408498 297978 409118 298046
rect 408498 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 409118 297978
rect 408498 280350 409118 297922
rect 408498 280294 408594 280350
rect 408650 280294 408718 280350
rect 408774 280294 408842 280350
rect 408898 280294 408966 280350
rect 409022 280294 409118 280350
rect 408498 280226 409118 280294
rect 408498 280170 408594 280226
rect 408650 280170 408718 280226
rect 408774 280170 408842 280226
rect 408898 280170 408966 280226
rect 409022 280170 409118 280226
rect 408498 280102 409118 280170
rect 408498 280046 408594 280102
rect 408650 280046 408718 280102
rect 408774 280046 408842 280102
rect 408898 280046 408966 280102
rect 409022 280046 409118 280102
rect 408498 279978 409118 280046
rect 408498 279922 408594 279978
rect 408650 279922 408718 279978
rect 408774 279922 408842 279978
rect 408898 279922 408966 279978
rect 409022 279922 409118 279978
rect 408498 262350 409118 279922
rect 408498 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 409118 262350
rect 408498 262226 409118 262294
rect 408498 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 409118 262226
rect 408498 262102 409118 262170
rect 408498 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 409118 262102
rect 408498 261978 409118 262046
rect 408498 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 409118 261978
rect 408498 244350 409118 261922
rect 435498 400350 436118 402722
rect 435498 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 436118 400350
rect 435498 400226 436118 400294
rect 435498 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 436118 400226
rect 435498 400102 436118 400170
rect 435498 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 436118 400102
rect 435498 399978 436118 400046
rect 435498 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 436118 399978
rect 435498 382350 436118 399922
rect 435498 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 436118 382350
rect 435498 382226 436118 382294
rect 435498 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 436118 382226
rect 435498 382102 436118 382170
rect 435498 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 436118 382102
rect 435498 381978 436118 382046
rect 435498 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 436118 381978
rect 435498 364350 436118 381922
rect 435498 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 436118 364350
rect 435498 364226 436118 364294
rect 435498 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 436118 364226
rect 435498 364102 436118 364170
rect 435498 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 436118 364102
rect 435498 363978 436118 364046
rect 435498 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 436118 363978
rect 435498 346350 436118 363922
rect 435498 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 436118 346350
rect 435498 346226 436118 346294
rect 435498 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 436118 346226
rect 435498 346102 436118 346170
rect 435498 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 436118 346102
rect 435498 345978 436118 346046
rect 435498 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 436118 345978
rect 435498 328350 436118 345922
rect 435498 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 436118 328350
rect 435498 328226 436118 328294
rect 435498 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 436118 328226
rect 435498 328102 436118 328170
rect 435498 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 436118 328102
rect 435498 327978 436118 328046
rect 435498 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 436118 327978
rect 435498 310350 436118 327922
rect 435498 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 436118 310350
rect 435498 310226 436118 310294
rect 435498 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 436118 310226
rect 435498 310102 436118 310170
rect 435498 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 436118 310102
rect 435498 309978 436118 310046
rect 435498 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 436118 309978
rect 435498 292350 436118 309922
rect 435498 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 436118 292350
rect 435498 292226 436118 292294
rect 435498 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 436118 292226
rect 435498 292102 436118 292170
rect 435498 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 436118 292102
rect 435498 291978 436118 292046
rect 435498 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 436118 291978
rect 435498 274350 436118 291922
rect 435498 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 436118 274350
rect 435498 274226 436118 274294
rect 435498 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 436118 274226
rect 435498 274102 436118 274170
rect 435498 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 436118 274102
rect 435498 273978 436118 274046
rect 435498 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 436118 273978
rect 408498 244294 408594 244350
rect 408650 244294 408718 244350
rect 408774 244294 408842 244350
rect 408898 244294 408966 244350
rect 409022 244294 409118 244350
rect 408498 244226 409118 244294
rect 408498 244170 408594 244226
rect 408650 244170 408718 244226
rect 408774 244170 408842 244226
rect 408898 244170 408966 244226
rect 409022 244170 409118 244226
rect 408498 244102 409118 244170
rect 408498 244046 408594 244102
rect 408650 244046 408718 244102
rect 408774 244046 408842 244102
rect 408898 244046 408966 244102
rect 409022 244046 409118 244102
rect 408498 243978 409118 244046
rect 408498 243922 408594 243978
rect 408650 243922 408718 243978
rect 408774 243922 408842 243978
rect 408898 243922 408966 243978
rect 409022 243922 409118 243978
rect 408498 226350 409118 243922
rect 408498 226294 408594 226350
rect 408650 226294 408718 226350
rect 408774 226294 408842 226350
rect 408898 226294 408966 226350
rect 409022 226294 409118 226350
rect 408498 226226 409118 226294
rect 408498 226170 408594 226226
rect 408650 226170 408718 226226
rect 408774 226170 408842 226226
rect 408898 226170 408966 226226
rect 409022 226170 409118 226226
rect 408498 226102 409118 226170
rect 408498 226046 408594 226102
rect 408650 226046 408718 226102
rect 408774 226046 408842 226102
rect 408898 226046 408966 226102
rect 409022 226046 409118 226102
rect 408498 225978 409118 226046
rect 408498 225922 408594 225978
rect 408650 225922 408718 225978
rect 408774 225922 408842 225978
rect 408898 225922 408966 225978
rect 409022 225922 409118 225978
rect 408498 208350 409118 225922
rect 408498 208294 408594 208350
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208294 409118 208350
rect 408498 208226 409118 208294
rect 408498 208170 408594 208226
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208170 409118 208226
rect 408498 208102 409118 208170
rect 408498 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 409118 208102
rect 408498 207978 409118 208046
rect 408498 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 409118 207978
rect 408498 190350 409118 207922
rect 408498 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 409118 190350
rect 408498 190226 409118 190294
rect 408498 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 409118 190226
rect 408498 190102 409118 190170
rect 408498 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 409118 190102
rect 408498 189978 409118 190046
rect 408498 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 409118 189978
rect 408498 172350 409118 189922
rect 408498 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 409118 172350
rect 408498 172226 409118 172294
rect 408498 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 409118 172226
rect 408498 172102 409118 172170
rect 408498 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 409118 172102
rect 408498 171978 409118 172046
rect 408498 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 409118 171978
rect 408498 154350 409118 171922
rect 408498 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 409118 154350
rect 408498 154226 409118 154294
rect 408498 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 409118 154226
rect 408498 154102 409118 154170
rect 408498 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 409118 154102
rect 408498 153978 409118 154046
rect 408498 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 409118 153978
rect 408498 136350 409118 153922
rect 412412 258804 412468 258814
rect 412412 142772 412468 258748
rect 412412 142706 412468 142716
rect 414092 258804 414148 258814
rect 414092 141204 414148 258748
rect 424396 258804 424452 258814
rect 424060 258468 424116 258478
rect 424060 255388 424116 258412
rect 424060 255332 424228 255388
rect 418348 142678 418404 142688
rect 418348 141958 418404 142622
rect 414092 141138 414148 141148
rect 414652 141204 414708 141214
rect 414652 141058 414708 141148
rect 418348 141204 418404 141902
rect 418348 141138 418404 141148
rect 414652 140992 414708 141002
rect 424172 139188 424228 255332
rect 424396 141876 424452 258748
rect 424396 141810 424452 141820
rect 433468 258692 433524 258702
rect 433468 140644 433524 258636
rect 434252 258580 434308 258590
rect 434140 258468 434196 258478
rect 434140 243628 434196 258412
rect 434252 255388 434308 258524
rect 434588 258468 434644 258478
rect 434252 255332 434420 255388
rect 433692 243572 434196 243628
rect 433692 142436 433748 243572
rect 433692 141988 433748 142380
rect 433692 141922 433748 141932
rect 434364 141764 434420 255332
rect 434364 141698 434420 141708
rect 434588 141764 434644 258412
rect 434588 141540 434644 141708
rect 434588 141474 434644 141484
rect 435498 256350 436118 273922
rect 435498 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 436118 256350
rect 435498 256226 436118 256294
rect 435498 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 436118 256226
rect 435498 256102 436118 256170
rect 435498 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 436118 256102
rect 435498 255978 436118 256046
rect 435498 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 436118 255978
rect 435498 238350 436118 255922
rect 435498 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 436118 238350
rect 435498 238226 436118 238294
rect 435498 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 436118 238226
rect 435498 238102 436118 238170
rect 435498 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 436118 238102
rect 435498 237978 436118 238046
rect 435498 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 436118 237978
rect 435498 220350 436118 237922
rect 435498 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 436118 220350
rect 435498 220226 436118 220294
rect 435498 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 436118 220226
rect 435498 220102 436118 220170
rect 435498 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 436118 220102
rect 435498 219978 436118 220046
rect 435498 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 436118 219978
rect 435498 202350 436118 219922
rect 435498 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 436118 202350
rect 435498 202226 436118 202294
rect 435498 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 436118 202226
rect 435498 202102 436118 202170
rect 435498 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 436118 202102
rect 435498 201978 436118 202046
rect 435498 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 436118 201978
rect 435498 184350 436118 201922
rect 435498 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 436118 184350
rect 435498 184226 436118 184294
rect 435498 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 436118 184226
rect 435498 184102 436118 184170
rect 435498 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 436118 184102
rect 435498 183978 436118 184046
rect 435498 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 436118 183978
rect 435498 166350 436118 183922
rect 435498 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 436118 166350
rect 435498 166226 436118 166294
rect 435498 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 436118 166226
rect 435498 166102 436118 166170
rect 435498 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 436118 166102
rect 435498 165978 436118 166046
rect 435498 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 436118 165978
rect 435498 148350 436118 165922
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 433468 140578 433524 140588
rect 424172 139122 424228 139132
rect 408498 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 409118 136350
rect 408498 136226 409118 136294
rect 408498 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 409118 136226
rect 408498 136102 409118 136170
rect 408498 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 409118 136102
rect 408498 135978 409118 136046
rect 408498 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 409118 135978
rect 408498 118350 409118 135922
rect 408498 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 409118 118350
rect 408498 118226 409118 118294
rect 408498 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 409118 118226
rect 408498 118102 409118 118170
rect 408498 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 409118 118102
rect 408498 117978 409118 118046
rect 408498 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 409118 117978
rect 408498 100350 409118 117922
rect 408498 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 409118 100350
rect 408498 100226 409118 100294
rect 408498 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 409118 100226
rect 408498 100102 409118 100170
rect 408498 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 409118 100102
rect 408498 99978 409118 100046
rect 408498 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 409118 99978
rect 408498 82350 409118 99922
rect 408498 82294 408594 82350
rect 408650 82294 408718 82350
rect 408774 82294 408842 82350
rect 408898 82294 408966 82350
rect 409022 82294 409118 82350
rect 408498 82226 409118 82294
rect 408498 82170 408594 82226
rect 408650 82170 408718 82226
rect 408774 82170 408842 82226
rect 408898 82170 408966 82226
rect 409022 82170 409118 82226
rect 408498 82102 409118 82170
rect 408498 82046 408594 82102
rect 408650 82046 408718 82102
rect 408774 82046 408842 82102
rect 408898 82046 408966 82102
rect 409022 82046 409118 82102
rect 408498 81978 409118 82046
rect 408498 81922 408594 81978
rect 408650 81922 408718 81978
rect 408774 81922 408842 81978
rect 408898 81922 408966 81978
rect 409022 81922 409118 81978
rect 408498 64350 409118 81922
rect 408498 64294 408594 64350
rect 408650 64294 408718 64350
rect 408774 64294 408842 64350
rect 408898 64294 408966 64350
rect 409022 64294 409118 64350
rect 408498 64226 409118 64294
rect 408498 64170 408594 64226
rect 408650 64170 408718 64226
rect 408774 64170 408842 64226
rect 408898 64170 408966 64226
rect 409022 64170 409118 64226
rect 408498 64102 409118 64170
rect 408498 64046 408594 64102
rect 408650 64046 408718 64102
rect 408774 64046 408842 64102
rect 408898 64046 408966 64102
rect 409022 64046 409118 64102
rect 408498 63978 409118 64046
rect 408498 63922 408594 63978
rect 408650 63922 408718 63978
rect 408774 63922 408842 63978
rect 408898 63922 408966 63978
rect 409022 63922 409118 63978
rect 408498 46350 409118 63922
rect 408498 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 409118 46350
rect 408498 46226 409118 46294
rect 408498 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 409118 46226
rect 408498 46102 409118 46170
rect 408498 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 409118 46102
rect 408498 45978 409118 46046
rect 408498 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 409118 45978
rect 408498 28350 409118 45922
rect 408498 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 409118 28350
rect 408498 28226 409118 28294
rect 408498 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 409118 28226
rect 408498 28102 409118 28170
rect 408498 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 409118 28102
rect 408498 27978 409118 28046
rect 408498 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 409118 27978
rect 408498 10350 409118 27922
rect 408498 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 409118 10350
rect 408498 10226 409118 10294
rect 408498 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 409118 10226
rect 408498 10102 409118 10170
rect 408498 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 409118 10102
rect 408498 9978 409118 10046
rect 408498 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 409118 9978
rect 408498 -1120 409118 9922
rect 408498 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 409118 -1120
rect 408498 -1244 409118 -1176
rect 408498 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 409118 -1244
rect 408498 -1368 409118 -1300
rect 408498 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 409118 -1368
rect 408498 -1492 409118 -1424
rect 408498 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 409118 -1492
rect 408498 -1644 409118 -1548
rect 435498 130350 436118 147922
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 435498 112350 436118 129922
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 435498 94350 436118 111922
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 435498 76350 436118 93922
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 435498 58350 436118 75922
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 435498 40350 436118 57922
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 435498 4350 436118 21922
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 435498 4102 436118 4170
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 388350 439838 402722
rect 439218 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 439838 388350
rect 439218 388226 439838 388294
rect 439218 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 439838 388226
rect 439218 388102 439838 388170
rect 439218 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 439838 388102
rect 439218 387978 439838 388046
rect 439218 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 439838 387978
rect 439218 370350 439838 387922
rect 449372 386148 449428 410284
rect 451052 387492 451108 411852
rect 456092 408772 456148 408782
rect 451052 387426 451108 387436
rect 452732 407204 452788 407214
rect 449372 386082 449428 386092
rect 452732 383460 452788 407148
rect 452732 383394 452788 383404
rect 454412 404068 454468 404078
rect 454412 380772 454468 404012
rect 456092 384804 456148 408716
rect 456092 384738 456148 384748
rect 454412 380706 454468 380716
rect 459452 379988 459508 557882
rect 466218 544350 466838 561922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 568350 470558 585922
rect 469938 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 470558 568350
rect 469938 568226 470558 568294
rect 469938 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 470558 568226
rect 469938 568102 470558 568170
rect 469938 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 470558 568102
rect 469938 567978 470558 568046
rect 469938 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 470558 567978
rect 469938 550350 470558 567922
rect 469938 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 470558 550350
rect 469938 550226 470558 550294
rect 469938 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 470558 550226
rect 469938 550102 470558 550170
rect 469938 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 470558 550102
rect 469938 549978 470558 550046
rect 469938 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 470558 549978
rect 468300 548996 468356 549006
rect 466218 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 466838 544350
rect 466218 544226 466838 544294
rect 466218 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 466838 544226
rect 466218 544102 466838 544170
rect 466218 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 466838 544102
rect 466218 543978 466838 544046
rect 466218 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 466838 543978
rect 466218 526350 466838 543922
rect 466218 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 466838 526350
rect 466218 526226 466838 526294
rect 466218 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 466838 526226
rect 466218 526102 466838 526170
rect 466218 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 466838 526102
rect 466218 525978 466838 526046
rect 466218 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 466838 525978
rect 466218 508350 466838 525922
rect 466218 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 466838 508350
rect 466218 508226 466838 508294
rect 466218 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 466838 508226
rect 466218 508102 466838 508170
rect 466218 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 466838 508102
rect 466218 507978 466838 508046
rect 466218 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 466838 507978
rect 466218 490350 466838 507922
rect 467628 548436 467684 548446
rect 467628 495572 467684 548380
rect 467628 495506 467684 495516
rect 468188 546868 468244 546878
rect 466218 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 466838 490350
rect 466218 490226 466838 490294
rect 466218 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 466838 490226
rect 466218 490102 466838 490170
rect 466218 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 466838 490102
rect 466218 489978 466838 490046
rect 466218 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 466838 489978
rect 466218 472350 466838 489922
rect 468188 483476 468244 546812
rect 468188 483410 468244 483420
rect 468300 477428 468356 548940
rect 468524 548884 468580 548894
rect 468524 514108 468580 548828
rect 469938 532350 470558 549922
rect 469938 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 470558 532350
rect 469938 532226 470558 532294
rect 469938 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 470558 532226
rect 469938 532102 470558 532170
rect 469938 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 470558 532102
rect 469938 531978 470558 532046
rect 469938 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 470558 531978
rect 469938 514350 470558 531922
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 496938 562350 497558 579922
rect 496938 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 497558 562350
rect 496938 562226 497558 562294
rect 496938 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 497558 562226
rect 496938 562102 497558 562170
rect 496938 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 497558 562102
rect 496938 561978 497558 562046
rect 496938 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 497558 561978
rect 496938 544350 497558 561922
rect 496938 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 497558 544350
rect 496938 544226 497558 544294
rect 496938 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 497558 544226
rect 496938 544102 497558 544170
rect 496938 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 497558 544102
rect 496938 543978 497558 544046
rect 496938 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 497558 543978
rect 496938 526432 497558 543922
rect 474448 526350 474768 526384
rect 474448 526294 474518 526350
rect 474574 526294 474642 526350
rect 474698 526294 474768 526350
rect 474448 526226 474768 526294
rect 496938 526376 497034 526432
rect 497090 526376 497158 526432
rect 497214 526376 497282 526432
rect 497338 526376 497406 526432
rect 497462 526376 497558 526432
rect 496938 526308 497558 526376
rect 496938 526252 497034 526308
rect 497090 526252 497158 526308
rect 497214 526252 497282 526308
rect 497338 526252 497406 526308
rect 497462 526252 497558 526308
rect 496938 526238 497558 526252
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 568350 501278 585922
rect 500658 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 501278 568350
rect 500658 568226 501278 568294
rect 500658 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 501278 568226
rect 500658 568102 501278 568170
rect 500658 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 501278 568102
rect 500658 567978 501278 568046
rect 500658 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 501278 567978
rect 500658 550350 501278 567922
rect 500658 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 501278 550350
rect 500658 550226 501278 550294
rect 500658 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 501278 550226
rect 500658 550102 501278 550170
rect 500658 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 501278 550102
rect 500658 549978 501278 550046
rect 500658 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 501278 549978
rect 500658 532350 501278 549922
rect 500658 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 501278 532350
rect 500658 532226 501278 532294
rect 500658 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 501278 532226
rect 500658 532102 501278 532170
rect 500658 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 501278 532102
rect 500658 531978 501278 532046
rect 500658 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 501278 531978
rect 500658 526238 501278 531922
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 527658 562350 528278 579922
rect 527658 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 528278 562350
rect 527658 562226 528278 562294
rect 527658 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 528278 562226
rect 527658 562102 528278 562170
rect 527658 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 528278 562102
rect 527658 561978 528278 562046
rect 527658 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 528278 561978
rect 527658 544350 528278 561922
rect 527658 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 528278 544350
rect 527658 544226 528278 544294
rect 527658 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 528278 544226
rect 527658 544102 528278 544170
rect 527658 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 528278 544102
rect 527658 543978 528278 544046
rect 527658 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 528278 543978
rect 527658 526432 528278 543922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 568350 531998 585922
rect 531378 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 531998 568350
rect 531378 568226 531998 568294
rect 531378 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 531998 568226
rect 531378 568102 531998 568170
rect 531378 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 531998 568102
rect 531378 567978 531998 568046
rect 531378 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 531998 567978
rect 531378 550350 531998 567922
rect 531378 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 531998 550350
rect 531378 550226 531998 550294
rect 531378 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 531998 550226
rect 531378 550102 531998 550170
rect 531378 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 531998 550102
rect 531378 549978 531998 550046
rect 531378 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 531998 549978
rect 529340 534324 529396 534334
rect 529340 533428 529396 534268
rect 529340 533362 529396 533372
rect 505168 526350 505488 526384
rect 505168 526294 505238 526350
rect 505294 526294 505362 526350
rect 505418 526294 505488 526350
rect 474448 526170 474518 526226
rect 474574 526170 474642 526226
rect 474698 526170 474768 526226
rect 474448 526102 474768 526170
rect 474448 526046 474518 526102
rect 474574 526046 474642 526102
rect 474698 526046 474768 526102
rect 474448 525978 474768 526046
rect 474448 525922 474518 525978
rect 474574 525922 474642 525978
rect 474698 525922 474768 525978
rect 474448 525888 474768 525922
rect 505168 526226 505488 526294
rect 527658 526376 527754 526432
rect 527810 526376 527878 526432
rect 527934 526376 528002 526432
rect 528058 526376 528126 526432
rect 528182 526376 528278 526432
rect 527658 526308 528278 526376
rect 527658 526252 527754 526308
rect 527810 526252 527878 526308
rect 527934 526252 528002 526308
rect 528058 526252 528126 526308
rect 528182 526252 528278 526308
rect 527658 526238 528278 526252
rect 531378 532350 531998 549922
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 558378 580350 558998 596784
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 556220 546418 556276 546428
rect 556108 546238 556164 546248
rect 531378 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 531998 532350
rect 531378 532226 531998 532294
rect 531378 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 531998 532226
rect 531378 532102 531998 532170
rect 531378 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 531998 532102
rect 531378 531978 531998 532046
rect 531378 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 531998 531978
rect 531378 526238 531998 531922
rect 548156 537796 548212 537806
rect 535888 526350 536208 526384
rect 535888 526294 535958 526350
rect 536014 526294 536082 526350
rect 536138 526294 536208 526350
rect 505168 526170 505238 526226
rect 505294 526170 505362 526226
rect 505418 526170 505488 526226
rect 505168 526102 505488 526170
rect 505168 526046 505238 526102
rect 505294 526046 505362 526102
rect 505418 526046 505488 526102
rect 505168 525978 505488 526046
rect 505168 525922 505238 525978
rect 505294 525922 505362 525978
rect 505418 525922 505488 525978
rect 505168 525888 505488 525922
rect 535888 526226 536208 526294
rect 535888 526170 535958 526226
rect 536014 526170 536082 526226
rect 536138 526170 536208 526226
rect 535888 526102 536208 526170
rect 535888 526046 535958 526102
rect 536014 526046 536082 526102
rect 536138 526046 536208 526102
rect 535888 525978 536208 526046
rect 535888 525922 535958 525978
rect 536014 525922 536082 525978
rect 536138 525922 536208 525978
rect 535888 525888 536208 525922
rect 469938 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 470558 514350
rect 469938 514226 470558 514294
rect 469938 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 470558 514226
rect 468524 514052 468692 514108
rect 468300 477362 468356 477372
rect 468636 489524 468692 514052
rect 466218 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 466838 472350
rect 466218 472226 466838 472294
rect 466218 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 466838 472226
rect 466218 472102 466838 472170
rect 466218 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 466838 472102
rect 466218 471978 466838 472046
rect 466218 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 466838 471978
rect 466218 454350 466838 471922
rect 466218 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 466838 454350
rect 466218 454226 466838 454294
rect 466218 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 466838 454226
rect 466218 454102 466838 454170
rect 466218 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 466838 454102
rect 466218 453978 466838 454046
rect 466218 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 466838 453978
rect 466218 436350 466838 453922
rect 466218 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 466838 436350
rect 466218 436226 466838 436294
rect 466218 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 466838 436226
rect 466218 436102 466838 436170
rect 466218 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 466838 436102
rect 466218 435978 466838 436046
rect 466218 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 466838 435978
rect 464604 430276 464660 430286
rect 459452 379922 459508 379932
rect 461132 429380 461188 429390
rect 439218 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 439838 370350
rect 439218 370226 439838 370294
rect 439218 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 439838 370226
rect 439218 370102 439838 370170
rect 439218 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 439838 370102
rect 439218 369978 439838 370046
rect 439218 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 439838 369978
rect 439218 352350 439838 369922
rect 451164 371458 451220 371468
rect 451052 364798 451108 364808
rect 439218 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 439838 352350
rect 439218 352226 439838 352294
rect 439218 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 439838 352226
rect 439218 352102 439838 352170
rect 439218 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 439838 352102
rect 439218 351978 439838 352046
rect 439218 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 439838 351978
rect 439218 334350 439838 351922
rect 449484 354538 449540 354548
rect 449372 343558 449428 343568
rect 439218 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 439838 334350
rect 439218 334226 439838 334294
rect 439218 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 439838 334226
rect 439218 334102 439838 334170
rect 439218 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 439838 334102
rect 439218 333978 439838 334046
rect 439218 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 439838 333978
rect 439218 316350 439838 333922
rect 439218 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 439838 316350
rect 439218 316226 439838 316294
rect 439218 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 439838 316226
rect 439218 316102 439838 316170
rect 439218 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 439838 316102
rect 439218 315978 439838 316046
rect 439218 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 439838 315978
rect 439218 298350 439838 315922
rect 439218 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 439838 298350
rect 439218 298226 439838 298294
rect 439218 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 439838 298226
rect 439218 298102 439838 298170
rect 439218 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 439838 298102
rect 439218 297978 439838 298046
rect 439218 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 439838 297978
rect 439218 280350 439838 297922
rect 439218 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 439838 280350
rect 439218 280226 439838 280294
rect 439218 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 439838 280226
rect 439218 280102 439838 280170
rect 439218 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 439838 280102
rect 439218 279978 439838 280046
rect 439218 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 439838 279978
rect 439218 262350 439838 279922
rect 439218 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 439838 262350
rect 439218 262226 439838 262294
rect 439218 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 439838 262226
rect 439218 262102 439838 262170
rect 439218 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 439838 262102
rect 439218 261978 439838 262046
rect 439218 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 439838 261978
rect 439218 244350 439838 261922
rect 447468 341938 447524 341948
rect 439218 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 439838 244350
rect 439218 244226 439838 244294
rect 439218 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 439838 244226
rect 439218 244102 439838 244170
rect 439218 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 439838 244102
rect 439218 243978 439838 244046
rect 439218 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 439838 243978
rect 439218 226350 439838 243922
rect 444668 258468 444724 258478
rect 444668 243628 444724 258412
rect 445340 258468 445396 258478
rect 445340 255388 445396 258412
rect 445340 255332 445620 255388
rect 439218 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 439838 226350
rect 439218 226226 439838 226294
rect 439218 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 439838 226226
rect 439218 226102 439838 226170
rect 439218 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 439838 226102
rect 439218 225978 439838 226046
rect 439218 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 439838 225978
rect 439218 208350 439838 225922
rect 439218 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 439838 208350
rect 439218 208226 439838 208294
rect 439218 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 439838 208226
rect 439218 208102 439838 208170
rect 439218 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 439838 208102
rect 439218 207978 439838 208046
rect 439218 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 439838 207978
rect 439218 190350 439838 207922
rect 439218 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 439838 190350
rect 439218 190226 439838 190294
rect 439218 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 439838 190226
rect 439218 190102 439838 190170
rect 439218 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 439838 190102
rect 439218 189978 439838 190046
rect 439218 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 439838 189978
rect 439218 172350 439838 189922
rect 439218 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 439838 172350
rect 439218 172226 439838 172294
rect 439218 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 439838 172226
rect 439218 172102 439838 172170
rect 439218 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 439838 172102
rect 439218 171978 439838 172046
rect 439218 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 439838 171978
rect 439218 154350 439838 171922
rect 444332 243572 444724 243628
rect 444332 161308 444388 243572
rect 444332 161252 444724 161308
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 444668 142498 444724 161252
rect 444668 141988 444724 142442
rect 444668 141922 444724 141932
rect 445564 142318 445620 255332
rect 446588 244350 447064 244384
rect 446588 244294 446612 244350
rect 446668 244294 446736 244350
rect 446792 244294 446860 244350
rect 446916 244294 446984 244350
rect 447040 244294 447064 244350
rect 446588 244226 447064 244294
rect 446588 244170 446612 244226
rect 446668 244170 446736 244226
rect 446792 244170 446860 244226
rect 446916 244170 446984 244226
rect 447040 244170 447064 244226
rect 446588 244102 447064 244170
rect 446588 244046 446612 244102
rect 446668 244046 446736 244102
rect 446792 244046 446860 244102
rect 446916 244046 446984 244102
rect 447040 244046 447064 244102
rect 446588 243978 447064 244046
rect 446588 243922 446612 243978
rect 446668 243922 446736 243978
rect 446792 243922 446860 243978
rect 446916 243922 446984 243978
rect 447040 243922 447064 243978
rect 446588 243888 447064 243922
rect 445788 238350 446264 238384
rect 445788 238294 445812 238350
rect 445868 238294 445936 238350
rect 445992 238294 446060 238350
rect 446116 238294 446184 238350
rect 446240 238294 446264 238350
rect 445788 238226 446264 238294
rect 445788 238170 445812 238226
rect 445868 238170 445936 238226
rect 445992 238170 446060 238226
rect 446116 238170 446184 238226
rect 446240 238170 446264 238226
rect 445788 238102 446264 238170
rect 445788 238046 445812 238102
rect 445868 238046 445936 238102
rect 445992 238046 446060 238102
rect 446116 238046 446184 238102
rect 446240 238046 446264 238102
rect 445788 237978 446264 238046
rect 445788 237922 445812 237978
rect 445868 237922 445936 237978
rect 445992 237922 446060 237978
rect 446116 237922 446184 237978
rect 446240 237922 446264 237978
rect 445788 237888 446264 237922
rect 446588 226350 447064 226384
rect 446588 226294 446612 226350
rect 446668 226294 446736 226350
rect 446792 226294 446860 226350
rect 446916 226294 446984 226350
rect 447040 226294 447064 226350
rect 446588 226226 447064 226294
rect 446588 226170 446612 226226
rect 446668 226170 446736 226226
rect 446792 226170 446860 226226
rect 446916 226170 446984 226226
rect 447040 226170 447064 226226
rect 446588 226102 447064 226170
rect 446588 226046 446612 226102
rect 446668 226046 446736 226102
rect 446792 226046 446860 226102
rect 446916 226046 446984 226102
rect 447040 226046 447064 226102
rect 446588 225978 447064 226046
rect 446588 225922 446612 225978
rect 446668 225922 446736 225978
rect 446792 225922 446860 225978
rect 446916 225922 446984 225978
rect 447040 225922 447064 225978
rect 446588 225888 447064 225922
rect 445788 220350 446264 220384
rect 445788 220294 445812 220350
rect 445868 220294 445936 220350
rect 445992 220294 446060 220350
rect 446116 220294 446184 220350
rect 446240 220294 446264 220350
rect 445788 220226 446264 220294
rect 445788 220170 445812 220226
rect 445868 220170 445936 220226
rect 445992 220170 446060 220226
rect 446116 220170 446184 220226
rect 446240 220170 446264 220226
rect 445788 220102 446264 220170
rect 445788 220046 445812 220102
rect 445868 220046 445936 220102
rect 445992 220046 446060 220102
rect 446116 220046 446184 220102
rect 446240 220046 446264 220102
rect 445788 219978 446264 220046
rect 445788 219922 445812 219978
rect 445868 219922 445936 219978
rect 445992 219922 446060 219978
rect 446116 219922 446184 219978
rect 446240 219922 446264 219978
rect 445788 219888 446264 219922
rect 446588 208350 447064 208384
rect 446588 208294 446612 208350
rect 446668 208294 446736 208350
rect 446792 208294 446860 208350
rect 446916 208294 446984 208350
rect 447040 208294 447064 208350
rect 446588 208226 447064 208294
rect 446588 208170 446612 208226
rect 446668 208170 446736 208226
rect 446792 208170 446860 208226
rect 446916 208170 446984 208226
rect 447040 208170 447064 208226
rect 446588 208102 447064 208170
rect 446588 208046 446612 208102
rect 446668 208046 446736 208102
rect 446792 208046 446860 208102
rect 446916 208046 446984 208102
rect 447040 208046 447064 208102
rect 446588 207978 447064 208046
rect 446588 207922 446612 207978
rect 446668 207922 446736 207978
rect 446792 207922 446860 207978
rect 446916 207922 446984 207978
rect 447040 207922 447064 207978
rect 446588 207888 447064 207922
rect 445788 202350 446264 202384
rect 445788 202294 445812 202350
rect 445868 202294 445936 202350
rect 445992 202294 446060 202350
rect 446116 202294 446184 202350
rect 446240 202294 446264 202350
rect 445788 202226 446264 202294
rect 445788 202170 445812 202226
rect 445868 202170 445936 202226
rect 445992 202170 446060 202226
rect 446116 202170 446184 202226
rect 446240 202170 446264 202226
rect 445788 202102 446264 202170
rect 445788 202046 445812 202102
rect 445868 202046 445936 202102
rect 445992 202046 446060 202102
rect 446116 202046 446184 202102
rect 446240 202046 446264 202102
rect 445788 201978 446264 202046
rect 445788 201922 445812 201978
rect 445868 201922 445936 201978
rect 445992 201922 446060 201978
rect 446116 201922 446184 201978
rect 446240 201922 446264 201978
rect 445788 201888 446264 201922
rect 446588 190350 447064 190384
rect 446588 190294 446612 190350
rect 446668 190294 446736 190350
rect 446792 190294 446860 190350
rect 446916 190294 446984 190350
rect 447040 190294 447064 190350
rect 446588 190226 447064 190294
rect 446588 190170 446612 190226
rect 446668 190170 446736 190226
rect 446792 190170 446860 190226
rect 446916 190170 446984 190226
rect 447040 190170 447064 190226
rect 446588 190102 447064 190170
rect 446588 190046 446612 190102
rect 446668 190046 446736 190102
rect 446792 190046 446860 190102
rect 446916 190046 446984 190102
rect 447040 190046 447064 190102
rect 446588 189978 447064 190046
rect 446588 189922 446612 189978
rect 446668 189922 446736 189978
rect 446792 189922 446860 189978
rect 446916 189922 446984 189978
rect 447040 189922 447064 189978
rect 446588 189888 447064 189922
rect 445788 184350 446264 184384
rect 445788 184294 445812 184350
rect 445868 184294 445936 184350
rect 445992 184294 446060 184350
rect 446116 184294 446184 184350
rect 446240 184294 446264 184350
rect 445788 184226 446264 184294
rect 445788 184170 445812 184226
rect 445868 184170 445936 184226
rect 445992 184170 446060 184226
rect 446116 184170 446184 184226
rect 446240 184170 446264 184226
rect 445788 184102 446264 184170
rect 445788 184046 445812 184102
rect 445868 184046 445936 184102
rect 445992 184046 446060 184102
rect 446116 184046 446184 184102
rect 446240 184046 446264 184102
rect 445788 183978 446264 184046
rect 445788 183922 445812 183978
rect 445868 183922 445936 183978
rect 445992 183922 446060 183978
rect 446116 183922 446184 183978
rect 446240 183922 446264 183978
rect 445788 183888 446264 183922
rect 446588 172350 447064 172384
rect 446588 172294 446612 172350
rect 446668 172294 446736 172350
rect 446792 172294 446860 172350
rect 446916 172294 446984 172350
rect 447040 172294 447064 172350
rect 446588 172226 447064 172294
rect 446588 172170 446612 172226
rect 446668 172170 446736 172226
rect 446792 172170 446860 172226
rect 446916 172170 446984 172226
rect 447040 172170 447064 172226
rect 446588 172102 447064 172170
rect 446588 172046 446612 172102
rect 446668 172046 446736 172102
rect 446792 172046 446860 172102
rect 446916 172046 446984 172102
rect 447040 172046 447064 172102
rect 446588 171978 447064 172046
rect 446588 171922 446612 171978
rect 446668 171922 446736 171978
rect 446792 171922 446860 171978
rect 446916 171922 446984 171978
rect 447040 171922 447064 171978
rect 446588 171888 447064 171922
rect 445788 166350 446264 166384
rect 445788 166294 445812 166350
rect 445868 166294 445936 166350
rect 445992 166294 446060 166350
rect 446116 166294 446184 166350
rect 446240 166294 446264 166350
rect 445788 166226 446264 166294
rect 445788 166170 445812 166226
rect 445868 166170 445936 166226
rect 445992 166170 446060 166226
rect 446116 166170 446184 166226
rect 446240 166170 446264 166226
rect 445788 166102 446264 166170
rect 445788 166046 445812 166102
rect 445868 166046 445936 166102
rect 445992 166046 446060 166102
rect 446116 166046 446184 166102
rect 446240 166046 446264 166102
rect 445788 165978 446264 166046
rect 445788 165922 445812 165978
rect 445868 165922 445936 165978
rect 445992 165922 446060 165978
rect 446116 165922 446184 165978
rect 446240 165922 446264 165978
rect 445788 165888 446264 165922
rect 445564 139076 445620 142262
rect 445564 139010 445620 139020
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 439218 118350 439838 135922
rect 445788 130350 446264 130384
rect 445788 130294 445812 130350
rect 445868 130294 445936 130350
rect 445992 130294 446060 130350
rect 446116 130294 446184 130350
rect 446240 130294 446264 130350
rect 445788 130226 446264 130294
rect 445788 130170 445812 130226
rect 445868 130170 445936 130226
rect 445992 130170 446060 130226
rect 446116 130170 446184 130226
rect 446240 130170 446264 130226
rect 445788 130102 446264 130170
rect 445788 130046 445812 130102
rect 445868 130046 445936 130102
rect 445992 130046 446060 130102
rect 446116 130046 446184 130102
rect 446240 130046 446264 130102
rect 445788 129978 446264 130046
rect 445788 129922 445812 129978
rect 445868 129922 445936 129978
rect 445992 129922 446060 129978
rect 446116 129922 446184 129978
rect 446240 129922 446264 129978
rect 445788 129888 446264 129922
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 439218 100350 439838 117922
rect 446588 118350 447064 118384
rect 446588 118294 446612 118350
rect 446668 118294 446736 118350
rect 446792 118294 446860 118350
rect 446916 118294 446984 118350
rect 447040 118294 447064 118350
rect 446588 118226 447064 118294
rect 446588 118170 446612 118226
rect 446668 118170 446736 118226
rect 446792 118170 446860 118226
rect 446916 118170 446984 118226
rect 447040 118170 447064 118226
rect 446588 118102 447064 118170
rect 446588 118046 446612 118102
rect 446668 118046 446736 118102
rect 446792 118046 446860 118102
rect 446916 118046 446984 118102
rect 447040 118046 447064 118102
rect 446588 117978 447064 118046
rect 446588 117922 446612 117978
rect 446668 117922 446736 117978
rect 446792 117922 446860 117978
rect 446916 117922 446984 117978
rect 447040 117922 447064 117978
rect 446588 117888 447064 117922
rect 445788 112350 446264 112384
rect 445788 112294 445812 112350
rect 445868 112294 445936 112350
rect 445992 112294 446060 112350
rect 446116 112294 446184 112350
rect 446240 112294 446264 112350
rect 445788 112226 446264 112294
rect 445788 112170 445812 112226
rect 445868 112170 445936 112226
rect 445992 112170 446060 112226
rect 446116 112170 446184 112226
rect 446240 112170 446264 112226
rect 445788 112102 446264 112170
rect 445788 112046 445812 112102
rect 445868 112046 445936 112102
rect 445992 112046 446060 112102
rect 446116 112046 446184 112102
rect 446240 112046 446264 112102
rect 445788 111978 446264 112046
rect 445788 111922 445812 111978
rect 445868 111922 445936 111978
rect 445992 111922 446060 111978
rect 446116 111922 446184 111978
rect 446240 111922 446264 111978
rect 445788 111888 446264 111922
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 439218 82350 439838 99922
rect 446588 100350 447064 100384
rect 446588 100294 446612 100350
rect 446668 100294 446736 100350
rect 446792 100294 446860 100350
rect 446916 100294 446984 100350
rect 447040 100294 447064 100350
rect 446588 100226 447064 100294
rect 446588 100170 446612 100226
rect 446668 100170 446736 100226
rect 446792 100170 446860 100226
rect 446916 100170 446984 100226
rect 447040 100170 447064 100226
rect 446588 100102 447064 100170
rect 446588 100046 446612 100102
rect 446668 100046 446736 100102
rect 446792 100046 446860 100102
rect 446916 100046 446984 100102
rect 447040 100046 447064 100102
rect 446588 99978 447064 100046
rect 446588 99922 446612 99978
rect 446668 99922 446736 99978
rect 446792 99922 446860 99978
rect 446916 99922 446984 99978
rect 447040 99922 447064 99978
rect 446588 99888 447064 99922
rect 445788 94350 446264 94384
rect 445788 94294 445812 94350
rect 445868 94294 445936 94350
rect 445992 94294 446060 94350
rect 446116 94294 446184 94350
rect 446240 94294 446264 94350
rect 445788 94226 446264 94294
rect 445788 94170 445812 94226
rect 445868 94170 445936 94226
rect 445992 94170 446060 94226
rect 446116 94170 446184 94226
rect 446240 94170 446264 94226
rect 445788 94102 446264 94170
rect 445788 94046 445812 94102
rect 445868 94046 445936 94102
rect 445992 94046 446060 94102
rect 446116 94046 446184 94102
rect 446240 94046 446264 94102
rect 445788 93978 446264 94046
rect 445788 93922 445812 93978
rect 445868 93922 445936 93978
rect 445992 93922 446060 93978
rect 446116 93922 446184 93978
rect 446240 93922 446264 93978
rect 445788 93888 446264 93922
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 439218 64350 439838 81922
rect 446588 82350 447064 82384
rect 446588 82294 446612 82350
rect 446668 82294 446736 82350
rect 446792 82294 446860 82350
rect 446916 82294 446984 82350
rect 447040 82294 447064 82350
rect 446588 82226 447064 82294
rect 446588 82170 446612 82226
rect 446668 82170 446736 82226
rect 446792 82170 446860 82226
rect 446916 82170 446984 82226
rect 447040 82170 447064 82226
rect 446588 82102 447064 82170
rect 446588 82046 446612 82102
rect 446668 82046 446736 82102
rect 446792 82046 446860 82102
rect 446916 82046 446984 82102
rect 447040 82046 447064 82102
rect 446588 81978 447064 82046
rect 446588 81922 446612 81978
rect 446668 81922 446736 81978
rect 446792 81922 446860 81978
rect 446916 81922 446984 81978
rect 447040 81922 447064 81978
rect 446588 81888 447064 81922
rect 445788 76350 446264 76384
rect 445788 76294 445812 76350
rect 445868 76294 445936 76350
rect 445992 76294 446060 76350
rect 446116 76294 446184 76350
rect 446240 76294 446264 76350
rect 445788 76226 446264 76294
rect 445788 76170 445812 76226
rect 445868 76170 445936 76226
rect 445992 76170 446060 76226
rect 446116 76170 446184 76226
rect 446240 76170 446264 76226
rect 445788 76102 446264 76170
rect 445788 76046 445812 76102
rect 445868 76046 445936 76102
rect 445992 76046 446060 76102
rect 446116 76046 446184 76102
rect 446240 76046 446264 76102
rect 445788 75978 446264 76046
rect 445788 75922 445812 75978
rect 445868 75922 445936 75978
rect 445992 75922 446060 75978
rect 446116 75922 446184 75978
rect 446240 75922 446264 75978
rect 445788 75888 446264 75922
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 439218 46350 439838 63922
rect 446588 64350 447064 64384
rect 446588 64294 446612 64350
rect 446668 64294 446736 64350
rect 446792 64294 446860 64350
rect 446916 64294 446984 64350
rect 447040 64294 447064 64350
rect 446588 64226 447064 64294
rect 446588 64170 446612 64226
rect 446668 64170 446736 64226
rect 446792 64170 446860 64226
rect 446916 64170 446984 64226
rect 447040 64170 447064 64226
rect 446588 64102 447064 64170
rect 446588 64046 446612 64102
rect 446668 64046 446736 64102
rect 446792 64046 446860 64102
rect 446916 64046 446984 64102
rect 447040 64046 447064 64102
rect 446588 63978 447064 64046
rect 446588 63922 446612 63978
rect 446668 63922 446736 63978
rect 446792 63922 446860 63978
rect 446916 63922 446984 63978
rect 447040 63922 447064 63978
rect 446588 63888 447064 63922
rect 445788 58350 446264 58384
rect 445788 58294 445812 58350
rect 445868 58294 445936 58350
rect 445992 58294 446060 58350
rect 446116 58294 446184 58350
rect 446240 58294 446264 58350
rect 445788 58226 446264 58294
rect 445788 58170 445812 58226
rect 445868 58170 445936 58226
rect 445992 58170 446060 58226
rect 446116 58170 446184 58226
rect 446240 58170 446264 58226
rect 445788 58102 446264 58170
rect 445788 58046 445812 58102
rect 445868 58046 445936 58102
rect 445992 58046 446060 58102
rect 446116 58046 446184 58102
rect 446240 58046 446264 58102
rect 445788 57978 446264 58046
rect 445788 57922 445812 57978
rect 445868 57922 445936 57978
rect 445992 57922 446060 57978
rect 446116 57922 446184 57978
rect 446240 57922 446264 57978
rect 445788 57888 446264 57922
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 439218 28350 439838 45922
rect 446588 46350 447064 46384
rect 446588 46294 446612 46350
rect 446668 46294 446736 46350
rect 446792 46294 446860 46350
rect 446916 46294 446984 46350
rect 447040 46294 447064 46350
rect 446588 46226 447064 46294
rect 446588 46170 446612 46226
rect 446668 46170 446736 46226
rect 446792 46170 446860 46226
rect 446916 46170 446984 46226
rect 447040 46170 447064 46226
rect 446588 46102 447064 46170
rect 446588 46046 446612 46102
rect 446668 46046 446736 46102
rect 446792 46046 446860 46102
rect 446916 46046 446984 46102
rect 447040 46046 447064 46102
rect 446588 45978 447064 46046
rect 446588 45922 446612 45978
rect 446668 45922 446736 45978
rect 446792 45922 446860 45978
rect 446916 45922 446984 45978
rect 447040 45922 447064 45978
rect 446588 45888 447064 45922
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 439218 10350 439838 27922
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 439218 -1120 439838 9922
rect 447468 4228 447524 341882
rect 449372 4340 449428 343502
rect 449484 39508 449540 354482
rect 449484 39442 449540 39452
rect 451052 24388 451108 364742
rect 451164 32788 451220 371402
rect 457884 368038 457940 368048
rect 454524 366418 454580 366428
rect 454412 364618 454468 364628
rect 451164 32722 451220 32732
rect 452732 358678 452788 358688
rect 451052 24322 451108 24332
rect 452732 4452 452788 358622
rect 452844 356338 452900 356348
rect 452844 6020 452900 356282
rect 452844 5954 452900 5964
rect 454412 5908 454468 364562
rect 454524 37940 454580 366362
rect 456204 361378 456260 361388
rect 454524 37874 454580 37884
rect 456092 353638 456148 353648
rect 454412 5842 454468 5852
rect 456092 4676 456148 353582
rect 456204 38052 456260 361322
rect 456204 37986 456260 37996
rect 457772 350218 457828 350228
rect 456092 4610 456148 4620
rect 457772 4564 457828 350162
rect 457884 34468 457940 367982
rect 461132 248518 461188 429324
rect 461132 248452 461188 248462
rect 464492 429268 464548 429278
rect 464492 206578 464548 429212
rect 464604 235198 464660 430220
rect 464604 235132 464660 235142
rect 466218 418350 466838 435922
rect 466218 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 466838 418350
rect 466218 418226 466838 418294
rect 466218 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 466838 418226
rect 466218 418102 466838 418170
rect 466218 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 466838 418102
rect 466218 417978 466838 418046
rect 466218 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 466838 417978
rect 466218 400350 466838 417922
rect 467852 471380 467908 471390
rect 467852 404398 467908 471324
rect 468636 450324 468692 489468
rect 468636 450258 468692 450268
rect 469938 514102 470558 514170
rect 469938 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 470558 514102
rect 469938 513978 470558 514046
rect 469938 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 470558 513978
rect 469938 496350 470558 513922
rect 489808 514350 490128 514384
rect 489808 514294 489878 514350
rect 489934 514294 490002 514350
rect 490058 514294 490128 514350
rect 489808 514226 490128 514294
rect 489808 514170 489878 514226
rect 489934 514170 490002 514226
rect 490058 514170 490128 514226
rect 489808 514102 490128 514170
rect 489808 514046 489878 514102
rect 489934 514046 490002 514102
rect 490058 514046 490128 514102
rect 489808 513978 490128 514046
rect 489808 513922 489878 513978
rect 489934 513922 490002 513978
rect 490058 513922 490128 513978
rect 489808 513888 490128 513922
rect 520528 514350 520848 514384
rect 520528 514294 520598 514350
rect 520654 514294 520722 514350
rect 520778 514294 520848 514350
rect 520528 514226 520848 514294
rect 520528 514170 520598 514226
rect 520654 514170 520722 514226
rect 520778 514170 520848 514226
rect 520528 514102 520848 514170
rect 520528 514046 520598 514102
rect 520654 514046 520722 514102
rect 520778 514046 520848 514102
rect 520528 513978 520848 514046
rect 520528 513922 520598 513978
rect 520654 513922 520722 513978
rect 520778 513922 520848 513978
rect 520528 513888 520848 513922
rect 474448 508350 474768 508384
rect 474448 508294 474518 508350
rect 474574 508294 474642 508350
rect 474698 508294 474768 508350
rect 474448 508226 474768 508294
rect 474448 508170 474518 508226
rect 474574 508170 474642 508226
rect 474698 508170 474768 508226
rect 474448 508102 474768 508170
rect 474448 508046 474518 508102
rect 474574 508046 474642 508102
rect 474698 508046 474768 508102
rect 474448 507978 474768 508046
rect 474448 507922 474518 507978
rect 474574 507922 474642 507978
rect 474698 507922 474768 507978
rect 474448 507888 474768 507922
rect 505168 508350 505488 508384
rect 505168 508294 505238 508350
rect 505294 508294 505362 508350
rect 505418 508294 505488 508350
rect 505168 508226 505488 508294
rect 505168 508170 505238 508226
rect 505294 508170 505362 508226
rect 505418 508170 505488 508226
rect 505168 508102 505488 508170
rect 505168 508046 505238 508102
rect 505294 508046 505362 508102
rect 505418 508046 505488 508102
rect 505168 507978 505488 508046
rect 505168 507922 505238 507978
rect 505294 507922 505362 507978
rect 505418 507922 505488 507978
rect 505168 507888 505488 507922
rect 535888 508350 536208 508384
rect 535888 508294 535958 508350
rect 536014 508294 536082 508350
rect 536138 508294 536208 508350
rect 535888 508226 536208 508294
rect 535888 508170 535958 508226
rect 536014 508170 536082 508226
rect 536138 508170 536208 508226
rect 535888 508102 536208 508170
rect 535888 508046 535958 508102
rect 536014 508046 536082 508102
rect 536138 508046 536208 508102
rect 535888 507978 536208 508046
rect 535888 507922 535958 507978
rect 536014 507922 536082 507978
rect 536138 507922 536208 507978
rect 535888 507888 536208 507922
rect 469938 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 470558 496350
rect 469938 496226 470558 496294
rect 469938 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 470558 496226
rect 469938 496102 470558 496170
rect 469938 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 470558 496102
rect 469938 495978 470558 496046
rect 469938 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 470558 495978
rect 469938 478350 470558 495922
rect 474908 499798 474964 499808
rect 474448 490350 474768 490384
rect 474448 490294 474518 490350
rect 474574 490294 474642 490350
rect 474698 490294 474768 490350
rect 474448 490226 474768 490294
rect 474448 490170 474518 490226
rect 474574 490170 474642 490226
rect 474698 490170 474768 490226
rect 474448 490102 474768 490170
rect 474448 490046 474518 490102
rect 474574 490046 474642 490102
rect 474698 490046 474768 490102
rect 474448 489978 474768 490046
rect 474448 489922 474518 489978
rect 474574 489922 474642 489978
rect 474698 489922 474768 489978
rect 474448 489888 474768 489922
rect 469938 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 470558 478350
rect 469938 478226 470558 478294
rect 469938 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 470558 478226
rect 469938 478102 470558 478170
rect 469938 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 470558 478102
rect 469938 477978 470558 478046
rect 469938 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 470558 477978
rect 469938 460350 470558 477922
rect 474448 472350 474768 472384
rect 474448 472294 474518 472350
rect 474574 472294 474642 472350
rect 474698 472294 474768 472350
rect 474448 472226 474768 472294
rect 474448 472170 474518 472226
rect 474574 472170 474642 472226
rect 474698 472170 474768 472226
rect 474448 472102 474768 472170
rect 474448 472046 474518 472102
rect 474574 472046 474642 472102
rect 474698 472046 474768 472102
rect 474448 471978 474768 472046
rect 474448 471922 474518 471978
rect 474574 471922 474642 471978
rect 474698 471922 474768 471978
rect 474448 471888 474768 471922
rect 469938 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 470558 460350
rect 469938 460226 470558 460294
rect 469938 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 470558 460226
rect 469938 460102 470558 460170
rect 469938 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 470558 460102
rect 469938 459978 470558 460046
rect 469938 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 470558 459978
rect 469938 442350 470558 459922
rect 474448 454350 474768 454384
rect 474448 454294 474518 454350
rect 474574 454294 474642 454350
rect 474698 454294 474768 454350
rect 474448 454226 474768 454294
rect 474448 454170 474518 454226
rect 474574 454170 474642 454226
rect 474698 454170 474768 454226
rect 474448 454102 474768 454170
rect 474448 454046 474518 454102
rect 474574 454046 474642 454102
rect 474698 454046 474768 454102
rect 474448 453978 474768 454046
rect 474448 453922 474518 453978
rect 474574 453922 474642 453978
rect 474698 453922 474768 453978
rect 474448 453888 474768 453922
rect 474908 450548 474964 499742
rect 489808 496350 490128 496384
rect 489808 496294 489878 496350
rect 489934 496294 490002 496350
rect 490058 496294 490128 496350
rect 489808 496226 490128 496294
rect 489808 496170 489878 496226
rect 489934 496170 490002 496226
rect 490058 496170 490128 496226
rect 489808 496102 490128 496170
rect 489808 496046 489878 496102
rect 489934 496046 490002 496102
rect 490058 496046 490128 496102
rect 489808 495978 490128 496046
rect 489808 495922 489878 495978
rect 489934 495922 490002 495978
rect 490058 495922 490128 495978
rect 489808 495888 490128 495922
rect 520528 496350 520848 496384
rect 520528 496294 520598 496350
rect 520654 496294 520722 496350
rect 520778 496294 520848 496350
rect 520528 496226 520848 496294
rect 520528 496170 520598 496226
rect 520654 496170 520722 496226
rect 520778 496170 520848 496226
rect 520528 496102 520848 496170
rect 520528 496046 520598 496102
rect 520654 496046 520722 496102
rect 520778 496046 520848 496102
rect 520528 495978 520848 496046
rect 520528 495922 520598 495978
rect 520654 495922 520722 495978
rect 520778 495922 520848 495978
rect 520528 495888 520848 495922
rect 505168 490350 505488 490384
rect 505168 490294 505238 490350
rect 505294 490294 505362 490350
rect 505418 490294 505488 490350
rect 505168 490226 505488 490294
rect 505168 490170 505238 490226
rect 505294 490170 505362 490226
rect 505418 490170 505488 490226
rect 505168 490102 505488 490170
rect 505168 490046 505238 490102
rect 505294 490046 505362 490102
rect 505418 490046 505488 490102
rect 505168 489978 505488 490046
rect 505168 489922 505238 489978
rect 505294 489922 505362 489978
rect 505418 489922 505488 489978
rect 505168 489888 505488 489922
rect 535888 490350 536208 490384
rect 535888 490294 535958 490350
rect 536014 490294 536082 490350
rect 536138 490294 536208 490350
rect 535888 490226 536208 490294
rect 535888 490170 535958 490226
rect 536014 490170 536082 490226
rect 536138 490170 536208 490226
rect 535888 490102 536208 490170
rect 535888 490046 535958 490102
rect 536014 490046 536082 490102
rect 536138 490046 536208 490102
rect 535888 489978 536208 490046
rect 535888 489922 535958 489978
rect 536014 489922 536082 489978
rect 536138 489922 536208 489978
rect 535888 489888 536208 489922
rect 489808 478350 490128 478384
rect 489808 478294 489878 478350
rect 489934 478294 490002 478350
rect 490058 478294 490128 478350
rect 489808 478226 490128 478294
rect 489808 478170 489878 478226
rect 489934 478170 490002 478226
rect 490058 478170 490128 478226
rect 489808 478102 490128 478170
rect 489808 478046 489878 478102
rect 489934 478046 490002 478102
rect 490058 478046 490128 478102
rect 489808 477978 490128 478046
rect 489808 477922 489878 477978
rect 489934 477922 490002 477978
rect 490058 477922 490128 477978
rect 489808 477888 490128 477922
rect 520528 478350 520848 478384
rect 520528 478294 520598 478350
rect 520654 478294 520722 478350
rect 520778 478294 520848 478350
rect 520528 478226 520848 478294
rect 520528 478170 520598 478226
rect 520654 478170 520722 478226
rect 520778 478170 520848 478226
rect 520528 478102 520848 478170
rect 520528 478046 520598 478102
rect 520654 478046 520722 478102
rect 520778 478046 520848 478102
rect 520528 477978 520848 478046
rect 520528 477922 520598 477978
rect 520654 477922 520722 477978
rect 520778 477922 520848 477978
rect 520528 477888 520848 477922
rect 505168 472350 505488 472384
rect 505168 472294 505238 472350
rect 505294 472294 505362 472350
rect 505418 472294 505488 472350
rect 505168 472226 505488 472294
rect 505168 472170 505238 472226
rect 505294 472170 505362 472226
rect 505418 472170 505488 472226
rect 505168 472102 505488 472170
rect 505168 472046 505238 472102
rect 505294 472046 505362 472102
rect 505418 472046 505488 472102
rect 505168 471978 505488 472046
rect 505168 471922 505238 471978
rect 505294 471922 505362 471978
rect 505418 471922 505488 471978
rect 505168 471888 505488 471922
rect 535888 472350 536208 472384
rect 535888 472294 535958 472350
rect 536014 472294 536082 472350
rect 536138 472294 536208 472350
rect 535888 472226 536208 472294
rect 535888 472170 535958 472226
rect 536014 472170 536082 472226
rect 536138 472170 536208 472226
rect 535888 472102 536208 472170
rect 535888 472046 535958 472102
rect 536014 472046 536082 472102
rect 536138 472046 536208 472102
rect 535888 471978 536208 472046
rect 535888 471922 535958 471978
rect 536014 471922 536082 471978
rect 536138 471922 536208 471978
rect 535888 471888 536208 471922
rect 489808 460350 490128 460384
rect 489808 460294 489878 460350
rect 489934 460294 490002 460350
rect 490058 460294 490128 460350
rect 489808 460226 490128 460294
rect 489808 460170 489878 460226
rect 489934 460170 490002 460226
rect 490058 460170 490128 460226
rect 489808 460102 490128 460170
rect 489808 460046 489878 460102
rect 489934 460046 490002 460102
rect 490058 460046 490128 460102
rect 489808 459978 490128 460046
rect 489808 459922 489878 459978
rect 489934 459922 490002 459978
rect 490058 459922 490128 459978
rect 489808 459888 490128 459922
rect 520528 460350 520848 460384
rect 520528 460294 520598 460350
rect 520654 460294 520722 460350
rect 520778 460294 520848 460350
rect 520528 460226 520848 460294
rect 520528 460170 520598 460226
rect 520654 460170 520722 460226
rect 520778 460170 520848 460226
rect 520528 460102 520848 460170
rect 520528 460046 520598 460102
rect 520654 460046 520722 460102
rect 520778 460046 520848 460102
rect 520528 459978 520848 460046
rect 520528 459922 520598 459978
rect 520654 459922 520722 459978
rect 520778 459922 520848 459978
rect 520528 459888 520848 459922
rect 505168 454350 505488 454384
rect 505168 454294 505238 454350
rect 505294 454294 505362 454350
rect 505418 454294 505488 454350
rect 505168 454226 505488 454294
rect 505168 454170 505238 454226
rect 505294 454170 505362 454226
rect 505418 454170 505488 454226
rect 505168 454102 505488 454170
rect 505168 454046 505238 454102
rect 505294 454046 505362 454102
rect 505418 454046 505488 454102
rect 505168 453978 505488 454046
rect 505168 453922 505238 453978
rect 505294 453922 505362 453978
rect 505418 453922 505488 453978
rect 505168 453888 505488 453922
rect 535888 454350 536208 454384
rect 535888 454294 535958 454350
rect 536014 454294 536082 454350
rect 536138 454294 536208 454350
rect 535888 454226 536208 454294
rect 535888 454170 535958 454226
rect 536014 454170 536082 454226
rect 536138 454170 536208 454226
rect 535888 454102 536208 454170
rect 535888 454046 535958 454102
rect 536014 454046 536082 454102
rect 536138 454046 536208 454102
rect 535888 453978 536208 454046
rect 535888 453922 535958 453978
rect 536014 453922 536082 453978
rect 536138 453922 536208 453978
rect 535888 453888 536208 453922
rect 481628 451444 481684 451454
rect 481404 451332 481460 451342
rect 481292 451108 481348 451118
rect 474908 450482 474964 450492
rect 478044 451018 478100 451028
rect 469938 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 470558 442350
rect 469938 442226 470558 442294
rect 469938 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 470558 442226
rect 469938 442102 470558 442170
rect 469938 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 470558 442102
rect 469938 441978 470558 442046
rect 469938 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 470558 441978
rect 469938 424350 470558 441922
rect 469938 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 470558 424350
rect 469938 424226 470558 424294
rect 469938 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 470558 424226
rect 469938 424102 470558 424170
rect 469938 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 470558 424102
rect 469938 423978 470558 424046
rect 469938 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 470558 423978
rect 469938 406350 470558 423922
rect 469938 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 470558 406350
rect 469938 406226 470558 406294
rect 469938 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 470558 406226
rect 469938 406102 470558 406170
rect 469938 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 470558 406102
rect 469938 405978 470558 406046
rect 469938 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 470558 405978
rect 467852 404332 467908 404342
rect 468636 404398 468692 404408
rect 468636 403396 468692 404342
rect 468636 403330 468692 403340
rect 466218 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 466838 400350
rect 466218 400226 466838 400294
rect 466218 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 466838 400226
rect 466218 400102 466838 400170
rect 466218 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 466838 400102
rect 466218 399978 466838 400046
rect 466218 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 466838 399978
rect 466218 382350 466838 399922
rect 466218 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 466838 382350
rect 466218 382226 466838 382294
rect 466218 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 466838 382226
rect 466218 382102 466838 382170
rect 466218 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 466838 382102
rect 466218 381978 466838 382046
rect 466218 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 466838 381978
rect 466218 364350 466838 381922
rect 466218 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 466838 364350
rect 466218 364226 466838 364294
rect 466218 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 466838 364226
rect 466218 364102 466838 364170
rect 466218 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 466838 364102
rect 466218 363978 466838 364046
rect 466218 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 466838 363978
rect 466218 346350 466838 363922
rect 466218 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 466838 346350
rect 466218 346226 466838 346294
rect 466218 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 466838 346226
rect 466218 346102 466838 346170
rect 466218 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 466838 346102
rect 466218 345978 466838 346046
rect 466218 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 466838 345978
rect 466218 328350 466838 345922
rect 466218 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 466838 328350
rect 466218 328226 466838 328294
rect 466218 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 466838 328226
rect 466218 328102 466838 328170
rect 466218 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 466838 328102
rect 466218 327978 466838 328046
rect 466218 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 466838 327978
rect 466218 310350 466838 327922
rect 466218 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 466838 310350
rect 466218 310226 466838 310294
rect 466218 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 466838 310226
rect 466218 310102 466838 310170
rect 466218 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 466838 310102
rect 466218 309978 466838 310046
rect 466218 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 466838 309978
rect 466218 292350 466838 309922
rect 466218 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 466838 292350
rect 466218 292226 466838 292294
rect 466218 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 466838 292226
rect 466218 292102 466838 292170
rect 466218 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 466838 292102
rect 466218 291978 466838 292046
rect 466218 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 466838 291978
rect 466218 274350 466838 291922
rect 466218 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 466838 274350
rect 466218 274226 466838 274294
rect 466218 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 466838 274226
rect 466218 274102 466838 274170
rect 466218 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 466838 274102
rect 466218 273978 466838 274046
rect 466218 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 466838 273978
rect 466218 256350 466838 273922
rect 466218 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 466838 256350
rect 466218 256226 466838 256294
rect 466218 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 466838 256226
rect 466218 256102 466838 256170
rect 466218 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 466838 256102
rect 466218 255978 466838 256046
rect 466218 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255922 466838 255978
rect 466218 238350 466838 255922
rect 466218 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 466838 238350
rect 466218 238226 466838 238294
rect 466218 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 466838 238226
rect 466218 238102 466838 238170
rect 466218 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 466838 238102
rect 466218 237978 466838 238046
rect 466218 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 466838 237978
rect 464492 206512 464548 206522
rect 466218 220350 466838 237922
rect 466218 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 466838 220350
rect 466218 220226 466838 220294
rect 466218 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 466838 220226
rect 466218 220102 466838 220170
rect 466218 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 466838 220102
rect 466218 219978 466838 220046
rect 466218 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 466838 219978
rect 466218 202350 466838 219922
rect 466218 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 466838 202350
rect 466218 202226 466838 202294
rect 466218 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 466838 202226
rect 466218 202102 466838 202170
rect 466218 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 466838 202102
rect 466218 201978 466838 202046
rect 466218 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 466838 201978
rect 466218 184350 466838 201922
rect 466218 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 466838 184350
rect 466218 184226 466838 184294
rect 466218 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 466838 184226
rect 466218 184102 466838 184170
rect 466218 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 466838 184102
rect 466218 183978 466838 184046
rect 466218 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 466838 183978
rect 466218 166350 466838 183922
rect 466218 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 466838 166350
rect 466218 166226 466838 166294
rect 466218 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 466838 166226
rect 466218 166102 466838 166170
rect 466218 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 466838 166102
rect 466218 165978 466838 166046
rect 466218 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 466838 165978
rect 466218 148350 466838 165922
rect 466218 148294 466314 148350
rect 466370 148294 466438 148350
rect 466494 148294 466562 148350
rect 466618 148294 466686 148350
rect 466742 148294 466838 148350
rect 466218 148226 466838 148294
rect 466218 148170 466314 148226
rect 466370 148170 466438 148226
rect 466494 148170 466562 148226
rect 466618 148170 466686 148226
rect 466742 148170 466838 148226
rect 466218 148102 466838 148170
rect 466218 148046 466314 148102
rect 466370 148046 466438 148102
rect 466494 148046 466562 148102
rect 466618 148046 466686 148102
rect 466742 148046 466838 148102
rect 466218 147978 466838 148046
rect 466218 147922 466314 147978
rect 466370 147922 466438 147978
rect 466494 147922 466562 147978
rect 466618 147922 466686 147978
rect 466742 147922 466838 147978
rect 461106 130350 461582 130384
rect 461106 130294 461130 130350
rect 461186 130294 461254 130350
rect 461310 130294 461378 130350
rect 461434 130294 461502 130350
rect 461558 130294 461582 130350
rect 461106 130226 461582 130294
rect 461106 130170 461130 130226
rect 461186 130170 461254 130226
rect 461310 130170 461378 130226
rect 461434 130170 461502 130226
rect 461558 130170 461582 130226
rect 461106 130102 461582 130170
rect 461106 130046 461130 130102
rect 461186 130046 461254 130102
rect 461310 130046 461378 130102
rect 461434 130046 461502 130102
rect 461558 130046 461582 130102
rect 461106 129978 461582 130046
rect 461106 129922 461130 129978
rect 461186 129922 461254 129978
rect 461310 129922 461378 129978
rect 461434 129922 461502 129978
rect 461558 129922 461582 129978
rect 461106 129888 461582 129922
rect 466218 130350 466838 147922
rect 466218 130294 466314 130350
rect 466370 130294 466438 130350
rect 466494 130294 466562 130350
rect 466618 130294 466686 130350
rect 466742 130294 466838 130350
rect 466218 130226 466838 130294
rect 466218 130170 466314 130226
rect 466370 130170 466438 130226
rect 466494 130170 466562 130226
rect 466618 130170 466686 130226
rect 466742 130170 466838 130226
rect 466218 130102 466838 130170
rect 466218 130046 466314 130102
rect 466370 130046 466438 130102
rect 466494 130046 466562 130102
rect 466618 130046 466686 130102
rect 466742 130046 466838 130102
rect 466218 129978 466838 130046
rect 466218 129922 466314 129978
rect 466370 129922 466438 129978
rect 466494 129922 466562 129978
rect 466618 129922 466686 129978
rect 466742 129922 466838 129978
rect 461906 118350 462382 118384
rect 461906 118294 461930 118350
rect 461986 118294 462054 118350
rect 462110 118294 462178 118350
rect 462234 118294 462302 118350
rect 462358 118294 462382 118350
rect 461906 118226 462382 118294
rect 461906 118170 461930 118226
rect 461986 118170 462054 118226
rect 462110 118170 462178 118226
rect 462234 118170 462302 118226
rect 462358 118170 462382 118226
rect 461906 118102 462382 118170
rect 461906 118046 461930 118102
rect 461986 118046 462054 118102
rect 462110 118046 462178 118102
rect 462234 118046 462302 118102
rect 462358 118046 462382 118102
rect 461906 117978 462382 118046
rect 461906 117922 461930 117978
rect 461986 117922 462054 117978
rect 462110 117922 462178 117978
rect 462234 117922 462302 117978
rect 462358 117922 462382 117978
rect 461906 117888 462382 117922
rect 461106 112350 461582 112384
rect 461106 112294 461130 112350
rect 461186 112294 461254 112350
rect 461310 112294 461378 112350
rect 461434 112294 461502 112350
rect 461558 112294 461582 112350
rect 461106 112226 461582 112294
rect 461106 112170 461130 112226
rect 461186 112170 461254 112226
rect 461310 112170 461378 112226
rect 461434 112170 461502 112226
rect 461558 112170 461582 112226
rect 461106 112102 461582 112170
rect 461106 112046 461130 112102
rect 461186 112046 461254 112102
rect 461310 112046 461378 112102
rect 461434 112046 461502 112102
rect 461558 112046 461582 112102
rect 461106 111978 461582 112046
rect 461106 111922 461130 111978
rect 461186 111922 461254 111978
rect 461310 111922 461378 111978
rect 461434 111922 461502 111978
rect 461558 111922 461582 111978
rect 461106 111888 461582 111922
rect 466218 112350 466838 129922
rect 466218 112294 466314 112350
rect 466370 112294 466438 112350
rect 466494 112294 466562 112350
rect 466618 112294 466686 112350
rect 466742 112294 466838 112350
rect 466218 112226 466838 112294
rect 466218 112170 466314 112226
rect 466370 112170 466438 112226
rect 466494 112170 466562 112226
rect 466618 112170 466686 112226
rect 466742 112170 466838 112226
rect 466218 112102 466838 112170
rect 466218 112046 466314 112102
rect 466370 112046 466438 112102
rect 466494 112046 466562 112102
rect 466618 112046 466686 112102
rect 466742 112046 466838 112102
rect 466218 111978 466838 112046
rect 466218 111922 466314 111978
rect 466370 111922 466438 111978
rect 466494 111922 466562 111978
rect 466618 111922 466686 111978
rect 466742 111922 466838 111978
rect 461906 100350 462382 100384
rect 461906 100294 461930 100350
rect 461986 100294 462054 100350
rect 462110 100294 462178 100350
rect 462234 100294 462302 100350
rect 462358 100294 462382 100350
rect 461906 100226 462382 100294
rect 461906 100170 461930 100226
rect 461986 100170 462054 100226
rect 462110 100170 462178 100226
rect 462234 100170 462302 100226
rect 462358 100170 462382 100226
rect 461906 100102 462382 100170
rect 461906 100046 461930 100102
rect 461986 100046 462054 100102
rect 462110 100046 462178 100102
rect 462234 100046 462302 100102
rect 462358 100046 462382 100102
rect 461906 99978 462382 100046
rect 461906 99922 461930 99978
rect 461986 99922 462054 99978
rect 462110 99922 462178 99978
rect 462234 99922 462302 99978
rect 462358 99922 462382 99978
rect 461906 99888 462382 99922
rect 461106 94350 461582 94384
rect 461106 94294 461130 94350
rect 461186 94294 461254 94350
rect 461310 94294 461378 94350
rect 461434 94294 461502 94350
rect 461558 94294 461582 94350
rect 461106 94226 461582 94294
rect 461106 94170 461130 94226
rect 461186 94170 461254 94226
rect 461310 94170 461378 94226
rect 461434 94170 461502 94226
rect 461558 94170 461582 94226
rect 461106 94102 461582 94170
rect 461106 94046 461130 94102
rect 461186 94046 461254 94102
rect 461310 94046 461378 94102
rect 461434 94046 461502 94102
rect 461558 94046 461582 94102
rect 461106 93978 461582 94046
rect 461106 93922 461130 93978
rect 461186 93922 461254 93978
rect 461310 93922 461378 93978
rect 461434 93922 461502 93978
rect 461558 93922 461582 93978
rect 461106 93888 461582 93922
rect 466218 94350 466838 111922
rect 466218 94294 466314 94350
rect 466370 94294 466438 94350
rect 466494 94294 466562 94350
rect 466618 94294 466686 94350
rect 466742 94294 466838 94350
rect 466218 94226 466838 94294
rect 466218 94170 466314 94226
rect 466370 94170 466438 94226
rect 466494 94170 466562 94226
rect 466618 94170 466686 94226
rect 466742 94170 466838 94226
rect 466218 94102 466838 94170
rect 466218 94046 466314 94102
rect 466370 94046 466438 94102
rect 466494 94046 466562 94102
rect 466618 94046 466686 94102
rect 466742 94046 466838 94102
rect 466218 93978 466838 94046
rect 466218 93922 466314 93978
rect 466370 93922 466438 93978
rect 466494 93922 466562 93978
rect 466618 93922 466686 93978
rect 466742 93922 466838 93978
rect 461906 82350 462382 82384
rect 461906 82294 461930 82350
rect 461986 82294 462054 82350
rect 462110 82294 462178 82350
rect 462234 82294 462302 82350
rect 462358 82294 462382 82350
rect 461906 82226 462382 82294
rect 461906 82170 461930 82226
rect 461986 82170 462054 82226
rect 462110 82170 462178 82226
rect 462234 82170 462302 82226
rect 462358 82170 462382 82226
rect 461906 82102 462382 82170
rect 461906 82046 461930 82102
rect 461986 82046 462054 82102
rect 462110 82046 462178 82102
rect 462234 82046 462302 82102
rect 462358 82046 462382 82102
rect 461906 81978 462382 82046
rect 461906 81922 461930 81978
rect 461986 81922 462054 81978
rect 462110 81922 462178 81978
rect 462234 81922 462302 81978
rect 462358 81922 462382 81978
rect 461906 81888 462382 81922
rect 461106 76350 461582 76384
rect 461106 76294 461130 76350
rect 461186 76294 461254 76350
rect 461310 76294 461378 76350
rect 461434 76294 461502 76350
rect 461558 76294 461582 76350
rect 461106 76226 461582 76294
rect 461106 76170 461130 76226
rect 461186 76170 461254 76226
rect 461310 76170 461378 76226
rect 461434 76170 461502 76226
rect 461558 76170 461582 76226
rect 461106 76102 461582 76170
rect 461106 76046 461130 76102
rect 461186 76046 461254 76102
rect 461310 76046 461378 76102
rect 461434 76046 461502 76102
rect 461558 76046 461582 76102
rect 461106 75978 461582 76046
rect 461106 75922 461130 75978
rect 461186 75922 461254 75978
rect 461310 75922 461378 75978
rect 461434 75922 461502 75978
rect 461558 75922 461582 75978
rect 461106 75888 461582 75922
rect 466218 76350 466838 93922
rect 466218 76294 466314 76350
rect 466370 76294 466438 76350
rect 466494 76294 466562 76350
rect 466618 76294 466686 76350
rect 466742 76294 466838 76350
rect 466218 76226 466838 76294
rect 466218 76170 466314 76226
rect 466370 76170 466438 76226
rect 466494 76170 466562 76226
rect 466618 76170 466686 76226
rect 466742 76170 466838 76226
rect 466218 76102 466838 76170
rect 466218 76046 466314 76102
rect 466370 76046 466438 76102
rect 466494 76046 466562 76102
rect 466618 76046 466686 76102
rect 466742 76046 466838 76102
rect 466218 75978 466838 76046
rect 466218 75922 466314 75978
rect 466370 75922 466438 75978
rect 466494 75922 466562 75978
rect 466618 75922 466686 75978
rect 466742 75922 466838 75978
rect 461906 64350 462382 64384
rect 461906 64294 461930 64350
rect 461986 64294 462054 64350
rect 462110 64294 462178 64350
rect 462234 64294 462302 64350
rect 462358 64294 462382 64350
rect 461906 64226 462382 64294
rect 461906 64170 461930 64226
rect 461986 64170 462054 64226
rect 462110 64170 462178 64226
rect 462234 64170 462302 64226
rect 462358 64170 462382 64226
rect 461906 64102 462382 64170
rect 461906 64046 461930 64102
rect 461986 64046 462054 64102
rect 462110 64046 462178 64102
rect 462234 64046 462302 64102
rect 462358 64046 462382 64102
rect 461906 63978 462382 64046
rect 461906 63922 461930 63978
rect 461986 63922 462054 63978
rect 462110 63922 462178 63978
rect 462234 63922 462302 63978
rect 462358 63922 462382 63978
rect 461906 63888 462382 63922
rect 461106 58350 461582 58384
rect 461106 58294 461130 58350
rect 461186 58294 461254 58350
rect 461310 58294 461378 58350
rect 461434 58294 461502 58350
rect 461558 58294 461582 58350
rect 461106 58226 461582 58294
rect 461106 58170 461130 58226
rect 461186 58170 461254 58226
rect 461310 58170 461378 58226
rect 461434 58170 461502 58226
rect 461558 58170 461582 58226
rect 461106 58102 461582 58170
rect 461106 58046 461130 58102
rect 461186 58046 461254 58102
rect 461310 58046 461378 58102
rect 461434 58046 461502 58102
rect 461558 58046 461582 58102
rect 461106 57978 461582 58046
rect 461106 57922 461130 57978
rect 461186 57922 461254 57978
rect 461310 57922 461378 57978
rect 461434 57922 461502 57978
rect 461558 57922 461582 57978
rect 461106 57888 461582 57922
rect 466218 58350 466838 75922
rect 466218 58294 466314 58350
rect 466370 58294 466438 58350
rect 466494 58294 466562 58350
rect 466618 58294 466686 58350
rect 466742 58294 466838 58350
rect 466218 58226 466838 58294
rect 466218 58170 466314 58226
rect 466370 58170 466438 58226
rect 466494 58170 466562 58226
rect 466618 58170 466686 58226
rect 466742 58170 466838 58226
rect 466218 58102 466838 58170
rect 466218 58046 466314 58102
rect 466370 58046 466438 58102
rect 466494 58046 466562 58102
rect 466618 58046 466686 58102
rect 466742 58046 466838 58102
rect 466218 57978 466838 58046
rect 466218 57922 466314 57978
rect 466370 57922 466438 57978
rect 466494 57922 466562 57978
rect 466618 57922 466686 57978
rect 466742 57922 466838 57978
rect 461906 46350 462382 46384
rect 461906 46294 461930 46350
rect 461986 46294 462054 46350
rect 462110 46294 462178 46350
rect 462234 46294 462302 46350
rect 462358 46294 462382 46350
rect 461906 46226 462382 46294
rect 461906 46170 461930 46226
rect 461986 46170 462054 46226
rect 462110 46170 462178 46226
rect 462234 46170 462302 46226
rect 462358 46170 462382 46226
rect 461906 46102 462382 46170
rect 461906 46046 461930 46102
rect 461986 46046 462054 46102
rect 462110 46046 462178 46102
rect 462234 46046 462302 46102
rect 462358 46046 462382 46102
rect 461906 45978 462382 46046
rect 461906 45922 461930 45978
rect 461986 45922 462054 45978
rect 462110 45922 462178 45978
rect 462234 45922 462302 45978
rect 462358 45922 462382 45978
rect 461906 45888 462382 45922
rect 457884 34402 457940 34412
rect 466218 40350 466838 57922
rect 466218 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 466838 40350
rect 466218 40226 466838 40294
rect 466218 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 466838 40226
rect 466218 40102 466838 40170
rect 466218 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 466838 40102
rect 466218 39978 466838 40046
rect 466218 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 466838 39978
rect 457772 4498 457828 4508
rect 466218 22350 466838 39922
rect 466218 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 466838 22350
rect 466218 22226 466838 22294
rect 466218 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 466838 22226
rect 466218 22102 466838 22170
rect 466218 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 466838 22102
rect 466218 21978 466838 22046
rect 466218 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 466838 21978
rect 452732 4386 452788 4396
rect 449372 4274 449428 4284
rect 466218 4350 466838 21922
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 447468 4162 447524 4172
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 388350 470558 405922
rect 474572 432292 474628 432302
rect 469938 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388294 470558 388350
rect 469938 388226 470558 388294
rect 469938 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 470558 388226
rect 469938 388102 470558 388170
rect 469938 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 470558 388102
rect 469938 387978 470558 388046
rect 469938 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 470558 387978
rect 469938 370350 470558 387922
rect 472892 402500 472948 402510
rect 472892 384020 472948 402444
rect 472892 383954 472948 383964
rect 469938 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 470558 370350
rect 469938 370226 470558 370294
rect 469938 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 470558 370226
rect 469938 370102 470558 370170
rect 469938 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 470558 370102
rect 469938 369978 470558 370046
rect 469938 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 470558 369978
rect 469938 352350 470558 369922
rect 469938 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 470558 352350
rect 469938 352226 470558 352294
rect 469938 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 470558 352226
rect 469938 352102 470558 352170
rect 469938 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 470558 352102
rect 469938 351978 470558 352046
rect 469938 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 470558 351978
rect 469938 334350 470558 351922
rect 469938 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 470558 334350
rect 469938 334226 470558 334294
rect 469938 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 470558 334226
rect 469938 334102 470558 334170
rect 469938 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 470558 334102
rect 469938 333978 470558 334046
rect 469938 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 470558 333978
rect 469938 316350 470558 333922
rect 469938 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 470558 316350
rect 469938 316226 470558 316294
rect 469938 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 470558 316226
rect 469938 316102 470558 316170
rect 469938 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 470558 316102
rect 469938 315978 470558 316046
rect 469938 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 470558 315978
rect 469938 298350 470558 315922
rect 469938 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 470558 298350
rect 469938 298226 470558 298294
rect 469938 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 470558 298226
rect 469938 298102 470558 298170
rect 469938 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 470558 298102
rect 469938 297978 470558 298046
rect 469938 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 470558 297978
rect 469938 280350 470558 297922
rect 472892 320516 472948 320526
rect 472892 280420 472948 320460
rect 473116 319620 473172 319630
rect 473116 280532 473172 319564
rect 474572 300538 474628 432236
rect 477932 431938 477988 431948
rect 474796 405636 474852 405646
rect 474684 400932 474740 400942
rect 474684 380660 474740 400876
rect 474796 390628 474852 405580
rect 474796 390562 474852 390572
rect 474684 380594 474740 380604
rect 475692 340318 475748 340328
rect 475468 339238 475524 339248
rect 475468 338436 475524 339182
rect 475468 338370 475524 338380
rect 475468 337618 475524 337628
rect 475468 337540 475524 337562
rect 475468 337474 475524 337484
rect 475580 337438 475636 337448
rect 475580 336644 475636 337382
rect 475580 336578 475636 336588
rect 475468 335998 475524 336008
rect 475468 335748 475524 335942
rect 475468 335682 475524 335692
rect 475468 333658 475524 333668
rect 475468 333060 475524 333602
rect 475468 332994 475524 333004
rect 475468 332578 475524 332588
rect 475468 332164 475524 332522
rect 475468 332098 475524 332108
rect 475580 332398 475636 332408
rect 475580 331268 475636 332342
rect 475580 331202 475636 331212
rect 475468 330958 475524 330968
rect 475468 330372 475524 330902
rect 475468 330306 475524 330316
rect 475692 329476 475748 340262
rect 475692 329410 475748 329420
rect 476252 340138 476308 340148
rect 476252 327684 476308 340082
rect 476252 327618 476308 327628
rect 475468 326788 475524 326798
rect 475468 326098 475524 326732
rect 475468 326032 475524 326042
rect 475468 321412 475524 321422
rect 475468 321058 475524 321356
rect 475468 320992 475524 321002
rect 475580 318724 475636 318734
rect 475468 317828 475524 317838
rect 475468 317734 475524 317762
rect 475580 317638 475636 318668
rect 475580 317572 475636 317582
rect 475468 315140 475524 315150
rect 475468 314218 475524 315084
rect 475468 314152 475524 314162
rect 475468 313348 475524 313358
rect 475468 312598 475524 313292
rect 475468 312532 475524 312542
rect 476588 311556 476644 311566
rect 476364 309764 476420 309774
rect 475468 308868 475524 308878
rect 475468 307558 475524 308812
rect 475468 307492 475524 307502
rect 476252 307972 476308 307982
rect 476140 305284 476196 305294
rect 476140 302428 476196 305228
rect 474572 300472 474628 300482
rect 476028 302372 476196 302428
rect 475468 289044 475524 289054
rect 475468 283618 475524 288988
rect 476028 288478 476084 302372
rect 476140 293972 476196 293982
rect 476140 290638 476196 293916
rect 476140 290572 476196 290582
rect 476028 288412 476084 288422
rect 475468 283552 475524 283562
rect 476252 281092 476308 307916
rect 476364 285418 476420 309708
rect 476364 285352 476420 285362
rect 476476 306180 476532 306190
rect 476252 281026 476308 281036
rect 476476 280756 476532 306124
rect 476588 287218 476644 311500
rect 476924 310660 476980 310670
rect 476700 307076 476756 307086
rect 476700 290458 476756 307020
rect 476700 290392 476756 290402
rect 476812 304388 476868 304398
rect 476588 287152 476644 287162
rect 476812 287038 476868 304332
rect 476924 293698 476980 310604
rect 476924 293632 476980 293642
rect 477036 303492 477092 303502
rect 476812 286972 476868 286982
rect 477036 286858 477092 303436
rect 477036 286792 477092 286802
rect 476476 280690 476532 280700
rect 473116 280466 473172 280476
rect 472892 280354 472948 280364
rect 469938 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 470558 280350
rect 469938 280226 470558 280294
rect 469938 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 470558 280226
rect 469938 280102 470558 280170
rect 469938 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 470558 280102
rect 469938 279978 470558 280046
rect 469938 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 470558 279978
rect 469938 262350 470558 279922
rect 477932 264740 477988 431882
rect 478044 399588 478100 450962
rect 478268 450660 478324 450670
rect 478044 399522 478100 399532
rect 478156 429492 478212 429502
rect 478156 398020 478212 429436
rect 478268 399476 478324 450604
rect 478492 450548 478548 450558
rect 478380 429940 478436 429950
rect 478380 401268 478436 429884
rect 478492 404578 478548 450492
rect 480508 450436 480564 450446
rect 479836 432478 479892 432488
rect 478492 404512 478548 404522
rect 479612 432298 479668 432308
rect 478380 401202 478436 401212
rect 478268 399410 478324 399420
rect 478156 397954 478212 397964
rect 478156 377524 478212 377534
rect 478156 288658 478212 377468
rect 478156 288592 478212 288602
rect 479612 269780 479668 432242
rect 479724 344596 479780 344606
rect 479724 295138 479780 344540
rect 479724 295072 479780 295082
rect 479836 283798 479892 432422
rect 480060 432118 480116 432128
rect 479948 344708 480004 344718
rect 479948 295318 480004 344652
rect 479948 295252 480004 295262
rect 480060 293878 480116 432062
rect 480508 401156 480564 450380
rect 480620 450324 480676 450334
rect 480620 420028 480676 450268
rect 480620 419972 480788 420028
rect 480620 405478 480676 405488
rect 480620 403172 480676 405422
rect 480620 403106 480676 403116
rect 480508 401090 480564 401100
rect 480508 400708 480564 400718
rect 480508 400438 480564 400652
rect 480732 400618 480788 419972
rect 481292 408268 481348 451052
rect 480620 400596 480788 400618
rect 480676 400562 480788 400596
rect 480844 408212 481348 408268
rect 480620 400530 480676 400540
rect 480844 400438 480900 408212
rect 481404 402958 481460 451276
rect 481516 451220 481572 451230
rect 481516 403138 481572 451164
rect 481628 405478 481684 451388
rect 526652 448532 526708 448542
rect 521612 447412 521668 447422
rect 512316 433378 512372 433388
rect 512316 432628 512372 433322
rect 512316 432562 512372 432572
rect 498876 432478 498932 432488
rect 481628 405412 481684 405422
rect 482972 432180 483028 432190
rect 481516 403072 481572 403082
rect 481404 402892 481460 402902
rect 480508 400382 480900 400438
rect 482972 398098 483028 432124
rect 498876 432180 498932 432422
rect 498876 432114 498932 432124
rect 502908 432298 502964 432308
rect 502908 432068 502964 432242
rect 502908 432002 502964 432012
rect 519036 432118 519092 432128
rect 519036 431956 519092 432062
rect 519036 431890 519092 431900
rect 483084 431844 483140 431854
rect 483084 402778 483140 431788
rect 499808 424350 500128 424384
rect 499808 424294 499878 424350
rect 499934 424294 500002 424350
rect 500058 424294 500128 424350
rect 499808 424226 500128 424294
rect 499808 424170 499878 424226
rect 499934 424170 500002 424226
rect 500058 424170 500128 424226
rect 499808 424102 500128 424170
rect 499808 424046 499878 424102
rect 499934 424046 500002 424102
rect 500058 424046 500128 424102
rect 499808 423978 500128 424046
rect 499808 423922 499878 423978
rect 499934 423922 500002 423978
rect 500058 423922 500128 423978
rect 499808 423888 500128 423922
rect 484448 418350 484768 418384
rect 484448 418294 484518 418350
rect 484574 418294 484642 418350
rect 484698 418294 484768 418350
rect 484448 418226 484768 418294
rect 484448 418170 484518 418226
rect 484574 418170 484642 418226
rect 484698 418170 484768 418226
rect 484448 418102 484768 418170
rect 484448 418046 484518 418102
rect 484574 418046 484642 418102
rect 484698 418046 484768 418102
rect 484448 417978 484768 418046
rect 484448 417922 484518 417978
rect 484574 417922 484642 417978
rect 484698 417922 484768 417978
rect 484448 417888 484768 417922
rect 515168 418350 515488 418384
rect 515168 418294 515238 418350
rect 515294 418294 515362 418350
rect 515418 418294 515488 418350
rect 515168 418226 515488 418294
rect 515168 418170 515238 418226
rect 515294 418170 515362 418226
rect 515418 418170 515488 418226
rect 515168 418102 515488 418170
rect 515168 418046 515238 418102
rect 515294 418046 515362 418102
rect 515418 418046 515488 418102
rect 515168 417978 515488 418046
rect 515168 417922 515238 417978
rect 515294 417922 515362 417978
rect 515418 417922 515488 417978
rect 515168 417888 515488 417922
rect 499808 406350 500128 406384
rect 499808 406294 499878 406350
rect 499934 406294 500002 406350
rect 500058 406294 500128 406350
rect 499808 406226 500128 406294
rect 499808 406170 499878 406226
rect 499934 406170 500002 406226
rect 500058 406170 500128 406226
rect 499808 406102 500128 406170
rect 499808 406046 499878 406102
rect 499934 406046 500002 406102
rect 500058 406046 500128 406102
rect 499808 405978 500128 406046
rect 499808 405922 499878 405978
rect 499934 405922 500002 405978
rect 500058 405922 500128 405978
rect 499808 405888 500128 405922
rect 483084 402712 483140 402722
rect 484448 400350 484768 400384
rect 484448 400294 484518 400350
rect 484574 400294 484642 400350
rect 484698 400294 484768 400350
rect 484448 400226 484768 400294
rect 484448 400170 484518 400226
rect 484574 400170 484642 400226
rect 484698 400170 484768 400226
rect 484448 400102 484768 400170
rect 484448 400046 484518 400102
rect 484574 400046 484642 400102
rect 484698 400046 484768 400102
rect 484448 399978 484768 400046
rect 484448 399922 484518 399978
rect 484574 399922 484642 399978
rect 484698 399922 484768 399978
rect 484448 399888 484768 399922
rect 515168 400350 515488 400384
rect 515168 400294 515238 400350
rect 515294 400294 515362 400350
rect 515418 400294 515488 400350
rect 515168 400226 515488 400294
rect 515168 400170 515238 400226
rect 515294 400170 515362 400226
rect 515418 400170 515488 400226
rect 515168 400102 515488 400170
rect 515168 400046 515238 400102
rect 515294 400046 515362 400102
rect 515418 400046 515488 400102
rect 515168 399978 515488 400046
rect 515168 399922 515238 399978
rect 515294 399922 515362 399978
rect 515418 399922 515488 399978
rect 515168 399888 515488 399922
rect 482972 398032 483028 398042
rect 499808 388350 500128 388384
rect 499808 388294 499878 388350
rect 499934 388294 500002 388350
rect 500058 388294 500128 388350
rect 499808 388226 500128 388294
rect 499808 388170 499878 388226
rect 499934 388170 500002 388226
rect 500058 388170 500128 388226
rect 499808 388102 500128 388170
rect 499808 388046 499878 388102
rect 499934 388046 500002 388102
rect 500058 388046 500128 388102
rect 499808 387978 500128 388046
rect 499808 387922 499878 387978
rect 499934 387922 500002 387978
rect 500058 387922 500128 387978
rect 499808 387888 500128 387922
rect 496938 382350 497558 387426
rect 496938 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 497558 382350
rect 496938 382226 497558 382294
rect 496938 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 497558 382226
rect 496938 382102 497558 382170
rect 496938 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 497558 382102
rect 496938 381978 497558 382046
rect 496938 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 497558 381978
rect 484764 381892 484820 381902
rect 484764 380772 484820 381836
rect 484764 380706 484820 380716
rect 494844 377972 494900 377982
rect 494844 377758 494900 377916
rect 494844 377692 494900 377702
rect 496938 364350 497558 381922
rect 498876 377972 498932 377982
rect 498876 377578 498932 377916
rect 498876 377512 498932 377522
rect 496938 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 497558 364350
rect 496938 364226 497558 364294
rect 496938 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 497558 364226
rect 496938 364102 497558 364170
rect 496938 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 497558 364102
rect 496938 363978 497558 364046
rect 496938 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 497558 363978
rect 495964 348598 496020 348608
rect 495964 344932 496020 348542
rect 495964 344866 496020 344876
rect 496938 346350 497558 363922
rect 500658 370350 501278 387426
rect 521052 377972 521108 377982
rect 521052 377872 521108 377882
rect 521612 377972 521668 447356
rect 523068 431938 523124 431948
rect 523068 431844 523124 431882
rect 523068 431778 523124 431788
rect 525868 388918 525924 388928
rect 525868 380436 525924 388862
rect 526652 388918 526708 448476
rect 526652 388852 526708 388862
rect 527658 436350 528278 453058
rect 527658 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 528278 436350
rect 527658 436226 528278 436294
rect 527658 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 528278 436226
rect 527658 436102 528278 436170
rect 527658 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 528278 436102
rect 527658 435978 528278 436046
rect 527658 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 528278 435978
rect 527658 418350 528278 435922
rect 527658 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 528278 418350
rect 527658 418226 528278 418294
rect 527658 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 528278 418226
rect 527658 418102 528278 418170
rect 527658 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 528278 418102
rect 527658 417978 528278 418046
rect 527658 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 528278 417978
rect 527658 400350 528278 417922
rect 527658 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 528278 400350
rect 527658 400226 528278 400294
rect 527658 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 528278 400226
rect 527658 400102 528278 400170
rect 527658 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 528278 400102
rect 527658 399978 528278 400046
rect 527658 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 528278 399978
rect 525868 380370 525924 380380
rect 527658 382350 528278 399922
rect 527658 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 528278 382350
rect 527658 382226 528278 382294
rect 527658 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 528278 382226
rect 527658 382102 528278 382170
rect 527658 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 528278 382102
rect 527658 381978 528278 382046
rect 527658 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 528278 381978
rect 500658 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 501278 370350
rect 500658 370226 501278 370294
rect 500658 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 501278 370226
rect 500658 370102 501278 370170
rect 500658 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 501278 370102
rect 500658 369978 501278 370046
rect 500658 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 501278 369978
rect 496938 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 497558 346350
rect 496938 346226 497558 346294
rect 496938 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 497558 346226
rect 496938 346102 497558 346170
rect 496938 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 497558 346102
rect 496938 345978 497558 346046
rect 496938 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 497558 345978
rect 480172 344484 480228 344494
rect 480172 298918 480228 344428
rect 496938 340062 497558 345922
rect 498988 360298 499044 360308
rect 498988 345380 499044 360242
rect 498988 345314 499044 345324
rect 500658 352350 501278 369922
rect 505708 373798 505764 373808
rect 500658 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 501278 352350
rect 500658 352226 501278 352294
rect 500658 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 501278 352226
rect 500658 352102 501278 352170
rect 500658 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 501278 352102
rect 500658 351978 501278 352046
rect 500658 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 501278 351978
rect 500658 340062 501278 351922
rect 502348 368758 502404 368768
rect 502348 345380 502404 368702
rect 502348 345314 502404 345324
rect 505708 345380 505764 373742
rect 521612 348628 521668 377916
rect 521612 348562 521668 348572
rect 527658 364350 528278 381922
rect 527658 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 528278 364350
rect 527658 364226 528278 364294
rect 527658 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 528278 364226
rect 527658 364102 528278 364170
rect 527658 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 528278 364102
rect 527658 363978 528278 364046
rect 527658 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 528278 363978
rect 527658 346350 528278 363922
rect 527658 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 528278 346350
rect 527658 346226 528278 346294
rect 527658 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 528278 346226
rect 527658 346102 528278 346170
rect 527658 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 528278 346102
rect 527658 345978 528278 346046
rect 527658 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 528278 345978
rect 519484 345718 519540 345728
rect 516124 345538 516180 345548
rect 505708 345314 505764 345324
rect 509404 345358 509460 345368
rect 509404 344484 509460 345302
rect 509404 344418 509460 344428
rect 512764 345178 512820 345188
rect 512764 344484 512820 345122
rect 512764 344418 512820 344428
rect 516124 344484 516180 345482
rect 516124 344418 516180 344428
rect 519484 344484 519540 345662
rect 519484 344418 519540 344428
rect 499808 334350 500128 334384
rect 499808 334294 499878 334350
rect 499934 334294 500002 334350
rect 500058 334294 500128 334350
rect 499808 334226 500128 334294
rect 499808 334170 499878 334226
rect 499934 334170 500002 334226
rect 500058 334170 500128 334226
rect 499808 334102 500128 334170
rect 499808 334046 499878 334102
rect 499934 334046 500002 334102
rect 500058 334046 500128 334102
rect 499808 333978 500128 334046
rect 499808 333922 499878 333978
rect 499934 333922 500002 333978
rect 500058 333922 500128 333978
rect 499808 333888 500128 333922
rect 484448 328350 484768 328384
rect 484448 328294 484518 328350
rect 484574 328294 484642 328350
rect 484698 328294 484768 328350
rect 484448 328226 484768 328294
rect 484448 328170 484518 328226
rect 484574 328170 484642 328226
rect 484698 328170 484768 328226
rect 484448 328102 484768 328170
rect 484448 328046 484518 328102
rect 484574 328046 484642 328102
rect 484698 328046 484768 328102
rect 484448 327978 484768 328046
rect 484448 327922 484518 327978
rect 484574 327922 484642 327978
rect 484698 327922 484768 327978
rect 484448 327888 484768 327922
rect 515168 328350 515488 328384
rect 515168 328294 515238 328350
rect 515294 328294 515362 328350
rect 515418 328294 515488 328350
rect 515168 328226 515488 328294
rect 515168 328170 515238 328226
rect 515294 328170 515362 328226
rect 515418 328170 515488 328226
rect 515168 328102 515488 328170
rect 515168 328046 515238 328102
rect 515294 328046 515362 328102
rect 515418 328046 515488 328102
rect 515168 327978 515488 328046
rect 515168 327922 515238 327978
rect 515294 327922 515362 327978
rect 515418 327922 515488 327978
rect 515168 327888 515488 327922
rect 527658 328350 528278 345922
rect 527658 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 528278 328350
rect 527658 328226 528278 328294
rect 527658 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 528278 328226
rect 527658 328102 528278 328170
rect 527658 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 528278 328102
rect 527658 327978 528278 328046
rect 527658 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 528278 327978
rect 499808 316350 500128 316384
rect 499808 316294 499878 316350
rect 499934 316294 500002 316350
rect 500058 316294 500128 316350
rect 499808 316226 500128 316294
rect 499808 316170 499878 316226
rect 499934 316170 500002 316226
rect 500058 316170 500128 316226
rect 499808 316102 500128 316170
rect 499808 316046 499878 316102
rect 499934 316046 500002 316102
rect 500058 316046 500128 316102
rect 499808 315978 500128 316046
rect 499808 315922 499878 315978
rect 499934 315922 500002 315978
rect 500058 315922 500128 315978
rect 499808 315888 500128 315922
rect 484448 310350 484768 310384
rect 484448 310294 484518 310350
rect 484574 310294 484642 310350
rect 484698 310294 484768 310350
rect 484448 310226 484768 310294
rect 484448 310170 484518 310226
rect 484574 310170 484642 310226
rect 484698 310170 484768 310226
rect 484448 310102 484768 310170
rect 484448 310046 484518 310102
rect 484574 310046 484642 310102
rect 484698 310046 484768 310102
rect 484448 309978 484768 310046
rect 484448 309922 484518 309978
rect 484574 309922 484642 309978
rect 484698 309922 484768 309978
rect 484448 309888 484768 309922
rect 515168 310350 515488 310384
rect 515168 310294 515238 310350
rect 515294 310294 515362 310350
rect 515418 310294 515488 310350
rect 515168 310226 515488 310294
rect 515168 310170 515238 310226
rect 515294 310170 515362 310226
rect 515418 310170 515488 310226
rect 515168 310102 515488 310170
rect 515168 310046 515238 310102
rect 515294 310046 515362 310102
rect 515418 310046 515488 310102
rect 515168 309978 515488 310046
rect 515168 309922 515238 309978
rect 515294 309922 515362 309978
rect 515418 309922 515488 309978
rect 515168 309888 515488 309922
rect 527658 310350 528278 327922
rect 527658 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 528278 310350
rect 527658 310226 528278 310294
rect 527658 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 528278 310226
rect 527658 310102 528278 310170
rect 527658 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 528278 310102
rect 527658 309978 528278 310046
rect 527658 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 528278 309978
rect 480172 298852 480228 298862
rect 480060 293812 480116 293822
rect 479836 283732 479892 283742
rect 496938 292350 497558 305970
rect 496938 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 497558 292350
rect 496938 292226 497558 292294
rect 496938 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 497558 292226
rect 496938 292102 497558 292170
rect 496938 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 497558 292102
rect 496938 291978 497558 292046
rect 496938 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 497558 291978
rect 479612 269714 479668 269724
rect 496938 274350 497558 291922
rect 496938 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 497558 274350
rect 496938 274226 497558 274294
rect 496938 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 497558 274226
rect 496938 274102 497558 274170
rect 496938 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 497558 274102
rect 496938 273978 497558 274046
rect 496938 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 497558 273978
rect 477932 264674 477988 264684
rect 469938 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 470558 262350
rect 469938 262226 470558 262294
rect 469938 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 470558 262226
rect 469938 262102 470558 262170
rect 469938 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 470558 262102
rect 469938 261978 470558 262046
rect 469938 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 470558 261978
rect 469938 244350 470558 261922
rect 496938 256350 497558 273922
rect 496938 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 497558 256350
rect 496938 256226 497558 256294
rect 496938 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 497558 256226
rect 496938 256102 497558 256170
rect 496938 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 497558 256102
rect 472708 256023 473184 256040
rect 472708 255967 472732 256023
rect 472788 255967 472856 256023
rect 472912 255967 472980 256023
rect 473036 255967 473104 256023
rect 473160 255967 473184 256023
rect 472708 255899 473184 255967
rect 472708 255843 472732 255899
rect 472788 255843 472856 255899
rect 472912 255843 472980 255899
rect 473036 255843 473104 255899
rect 473160 255843 473184 255899
rect 472708 255826 473184 255843
rect 496938 255978 497558 256046
rect 496938 255922 497034 255978
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 497558 255978
rect 469938 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 470558 244350
rect 469938 244226 470558 244294
rect 469938 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 470558 244226
rect 469938 244102 470558 244170
rect 469938 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 470558 244102
rect 469938 243978 470558 244046
rect 469938 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 470558 243978
rect 469938 226350 470558 243922
rect 471908 244350 472384 244384
rect 471908 244294 471932 244350
rect 471988 244294 472056 244350
rect 472112 244294 472180 244350
rect 472236 244294 472304 244350
rect 472360 244294 472384 244350
rect 471908 244226 472384 244294
rect 471908 244170 471932 244226
rect 471988 244170 472056 244226
rect 472112 244170 472180 244226
rect 472236 244170 472304 244226
rect 472360 244170 472384 244226
rect 471908 244102 472384 244170
rect 471908 244046 471932 244102
rect 471988 244046 472056 244102
rect 472112 244046 472180 244102
rect 472236 244046 472304 244102
rect 472360 244046 472384 244102
rect 471908 243978 472384 244046
rect 471908 243922 471932 243978
rect 471988 243922 472056 243978
rect 472112 243922 472180 243978
rect 472236 243922 472304 243978
rect 472360 243922 472384 243978
rect 471908 243888 472384 243922
rect 472708 238350 473184 238384
rect 472708 238294 472732 238350
rect 472788 238294 472856 238350
rect 472912 238294 472980 238350
rect 473036 238294 473104 238350
rect 473160 238294 473184 238350
rect 472708 238226 473184 238294
rect 472708 238170 472732 238226
rect 472788 238170 472856 238226
rect 472912 238170 472980 238226
rect 473036 238170 473104 238226
rect 473160 238170 473184 238226
rect 472708 238102 473184 238170
rect 472708 238046 472732 238102
rect 472788 238046 472856 238102
rect 472912 238046 472980 238102
rect 473036 238046 473104 238102
rect 473160 238046 473184 238102
rect 472708 237978 473184 238046
rect 472708 237922 472732 237978
rect 472788 237922 472856 237978
rect 472912 237922 472980 237978
rect 473036 237922 473104 237978
rect 473160 237922 473184 237978
rect 472708 237888 473184 237922
rect 496938 238350 497558 255922
rect 496938 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 497558 238350
rect 496938 238226 497558 238294
rect 496938 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 497558 238226
rect 496938 238102 497558 238170
rect 496938 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 497558 238102
rect 496938 237978 497558 238046
rect 496938 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 497558 237978
rect 469938 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 470558 226350
rect 469938 226226 470558 226294
rect 469938 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 470558 226226
rect 469938 226102 470558 226170
rect 469938 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 470558 226102
rect 469938 225978 470558 226046
rect 469938 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 470558 225978
rect 469938 208350 470558 225922
rect 471908 226350 472384 226384
rect 471908 226294 471932 226350
rect 471988 226294 472056 226350
rect 472112 226294 472180 226350
rect 472236 226294 472304 226350
rect 472360 226294 472384 226350
rect 471908 226226 472384 226294
rect 471908 226170 471932 226226
rect 471988 226170 472056 226226
rect 472112 226170 472180 226226
rect 472236 226170 472304 226226
rect 472360 226170 472384 226226
rect 471908 226102 472384 226170
rect 471908 226046 471932 226102
rect 471988 226046 472056 226102
rect 472112 226046 472180 226102
rect 472236 226046 472304 226102
rect 472360 226046 472384 226102
rect 471908 225978 472384 226046
rect 471908 225922 471932 225978
rect 471988 225922 472056 225978
rect 472112 225922 472180 225978
rect 472236 225922 472304 225978
rect 472360 225922 472384 225978
rect 471908 225888 472384 225922
rect 472708 220350 473184 220384
rect 472708 220294 472732 220350
rect 472788 220294 472856 220350
rect 472912 220294 472980 220350
rect 473036 220294 473104 220350
rect 473160 220294 473184 220350
rect 472708 220226 473184 220294
rect 472708 220170 472732 220226
rect 472788 220170 472856 220226
rect 472912 220170 472980 220226
rect 473036 220170 473104 220226
rect 473160 220170 473184 220226
rect 472708 220102 473184 220170
rect 472708 220046 472732 220102
rect 472788 220046 472856 220102
rect 472912 220046 472980 220102
rect 473036 220046 473104 220102
rect 473160 220046 473184 220102
rect 472708 219978 473184 220046
rect 472708 219922 472732 219978
rect 472788 219922 472856 219978
rect 472912 219922 472980 219978
rect 473036 219922 473104 219978
rect 473160 219922 473184 219978
rect 472708 219888 473184 219922
rect 496938 220350 497558 237922
rect 496938 220294 497034 220350
rect 497090 220294 497158 220350
rect 497214 220294 497282 220350
rect 497338 220294 497406 220350
rect 497462 220294 497558 220350
rect 496938 220226 497558 220294
rect 496938 220170 497034 220226
rect 497090 220170 497158 220226
rect 497214 220170 497282 220226
rect 497338 220170 497406 220226
rect 497462 220170 497558 220226
rect 496938 220102 497558 220170
rect 496938 220046 497034 220102
rect 497090 220046 497158 220102
rect 497214 220046 497282 220102
rect 497338 220046 497406 220102
rect 497462 220046 497558 220102
rect 496938 219978 497558 220046
rect 496938 219922 497034 219978
rect 497090 219922 497158 219978
rect 497214 219922 497282 219978
rect 497338 219922 497406 219978
rect 497462 219922 497558 219978
rect 469938 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 470558 208350
rect 469938 208226 470558 208294
rect 469938 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 470558 208226
rect 469938 208102 470558 208170
rect 469938 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 470558 208102
rect 469938 207978 470558 208046
rect 469938 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 470558 207978
rect 469938 190350 470558 207922
rect 471908 208350 472384 208384
rect 471908 208294 471932 208350
rect 471988 208294 472056 208350
rect 472112 208294 472180 208350
rect 472236 208294 472304 208350
rect 472360 208294 472384 208350
rect 471908 208226 472384 208294
rect 471908 208170 471932 208226
rect 471988 208170 472056 208226
rect 472112 208170 472180 208226
rect 472236 208170 472304 208226
rect 472360 208170 472384 208226
rect 471908 208102 472384 208170
rect 471908 208046 471932 208102
rect 471988 208046 472056 208102
rect 472112 208046 472180 208102
rect 472236 208046 472304 208102
rect 472360 208046 472384 208102
rect 471908 207978 472384 208046
rect 471908 207922 471932 207978
rect 471988 207922 472056 207978
rect 472112 207922 472180 207978
rect 472236 207922 472304 207978
rect 472360 207922 472384 207978
rect 471908 207888 472384 207922
rect 472708 202350 473184 202384
rect 472708 202294 472732 202350
rect 472788 202294 472856 202350
rect 472912 202294 472980 202350
rect 473036 202294 473104 202350
rect 473160 202294 473184 202350
rect 472708 202226 473184 202294
rect 472708 202170 472732 202226
rect 472788 202170 472856 202226
rect 472912 202170 472980 202226
rect 473036 202170 473104 202226
rect 473160 202170 473184 202226
rect 472708 202102 473184 202170
rect 472708 202046 472732 202102
rect 472788 202046 472856 202102
rect 472912 202046 472980 202102
rect 473036 202046 473104 202102
rect 473160 202046 473184 202102
rect 472708 201978 473184 202046
rect 472708 201922 472732 201978
rect 472788 201922 472856 201978
rect 472912 201922 472980 201978
rect 473036 201922 473104 201978
rect 473160 201922 473184 201978
rect 472708 201888 473184 201922
rect 496938 202350 497558 219922
rect 496938 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 497558 202350
rect 496938 202226 497558 202294
rect 496938 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 497558 202226
rect 496938 202102 497558 202170
rect 496938 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 497558 202102
rect 496938 201978 497558 202046
rect 496938 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 497558 201978
rect 469938 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 470558 190350
rect 469938 190226 470558 190294
rect 469938 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 470558 190226
rect 469938 190102 470558 190170
rect 469938 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 470558 190102
rect 469938 189978 470558 190046
rect 469938 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 470558 189978
rect 469938 172350 470558 189922
rect 471908 190350 472384 190384
rect 471908 190294 471932 190350
rect 471988 190294 472056 190350
rect 472112 190294 472180 190350
rect 472236 190294 472304 190350
rect 472360 190294 472384 190350
rect 471908 190226 472384 190294
rect 471908 190170 471932 190226
rect 471988 190170 472056 190226
rect 472112 190170 472180 190226
rect 472236 190170 472304 190226
rect 472360 190170 472384 190226
rect 471908 190102 472384 190170
rect 471908 190046 471932 190102
rect 471988 190046 472056 190102
rect 472112 190046 472180 190102
rect 472236 190046 472304 190102
rect 472360 190046 472384 190102
rect 471908 189978 472384 190046
rect 471908 189922 471932 189978
rect 471988 189922 472056 189978
rect 472112 189922 472180 189978
rect 472236 189922 472304 189978
rect 472360 189922 472384 189978
rect 471908 189888 472384 189922
rect 472708 184350 473184 184384
rect 472708 184294 472732 184350
rect 472788 184294 472856 184350
rect 472912 184294 472980 184350
rect 473036 184294 473104 184350
rect 473160 184294 473184 184350
rect 472708 184226 473184 184294
rect 472708 184170 472732 184226
rect 472788 184170 472856 184226
rect 472912 184170 472980 184226
rect 473036 184170 473104 184226
rect 473160 184170 473184 184226
rect 472708 184102 473184 184170
rect 472708 184046 472732 184102
rect 472788 184046 472856 184102
rect 472912 184046 472980 184102
rect 473036 184046 473104 184102
rect 473160 184046 473184 184102
rect 472708 183978 473184 184046
rect 472708 183922 472732 183978
rect 472788 183922 472856 183978
rect 472912 183922 472980 183978
rect 473036 183922 473104 183978
rect 473160 183922 473184 183978
rect 472708 183888 473184 183922
rect 496938 184350 497558 201922
rect 496938 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 497558 184350
rect 496938 184226 497558 184294
rect 496938 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 497558 184226
rect 496938 184102 497558 184170
rect 496938 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 497558 184102
rect 496938 183978 497558 184046
rect 496938 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 497558 183978
rect 469938 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 470558 172350
rect 469938 172226 470558 172294
rect 469938 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 470558 172226
rect 469938 172102 470558 172170
rect 469938 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 470558 172102
rect 469938 171978 470558 172046
rect 469938 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 470558 171978
rect 469938 154350 470558 171922
rect 471908 172350 472384 172384
rect 471908 172294 471932 172350
rect 471988 172294 472056 172350
rect 472112 172294 472180 172350
rect 472236 172294 472304 172350
rect 472360 172294 472384 172350
rect 471908 172226 472384 172294
rect 471908 172170 471932 172226
rect 471988 172170 472056 172226
rect 472112 172170 472180 172226
rect 472236 172170 472304 172226
rect 472360 172170 472384 172226
rect 471908 172102 472384 172170
rect 471908 172046 471932 172102
rect 471988 172046 472056 172102
rect 472112 172046 472180 172102
rect 472236 172046 472304 172102
rect 472360 172046 472384 172102
rect 471908 171978 472384 172046
rect 471908 171922 471932 171978
rect 471988 171922 472056 171978
rect 472112 171922 472180 171978
rect 472236 171922 472304 171978
rect 472360 171922 472384 171978
rect 471908 171888 472384 171922
rect 472708 166350 473184 166384
rect 472708 166294 472732 166350
rect 472788 166294 472856 166350
rect 472912 166294 472980 166350
rect 473036 166294 473104 166350
rect 473160 166294 473184 166350
rect 472708 166226 473184 166294
rect 472708 166170 472732 166226
rect 472788 166170 472856 166226
rect 472912 166170 472980 166226
rect 473036 166170 473104 166226
rect 473160 166170 473184 166226
rect 472708 166102 473184 166170
rect 472708 166046 472732 166102
rect 472788 166046 472856 166102
rect 472912 166046 472980 166102
rect 473036 166046 473104 166102
rect 473160 166046 473184 166102
rect 472708 165978 473184 166046
rect 472708 165922 472732 165978
rect 472788 165922 472856 165978
rect 472912 165922 472980 165978
rect 473036 165922 473104 165978
rect 473160 165922 473184 165978
rect 472708 165888 473184 165922
rect 496938 166350 497558 183922
rect 496938 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 497558 166350
rect 496938 166226 497558 166294
rect 496938 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 497558 166226
rect 496938 166102 497558 166170
rect 496938 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 497558 166102
rect 496938 165978 497558 166046
rect 496938 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 497558 165978
rect 469938 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 470558 154350
rect 469938 154226 470558 154294
rect 469938 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 470558 154226
rect 469938 154102 470558 154170
rect 469938 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 470558 154102
rect 469938 153978 470558 154046
rect 469938 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 470558 153978
rect 469938 136350 470558 153922
rect 474572 156324 474628 156334
rect 474572 142498 474628 156268
rect 474572 142432 474628 142442
rect 496938 148350 497558 165922
rect 496938 148294 497034 148350
rect 497090 148294 497158 148350
rect 497214 148294 497282 148350
rect 497338 148294 497406 148350
rect 497462 148294 497558 148350
rect 496938 148226 497558 148294
rect 496938 148170 497034 148226
rect 497090 148170 497158 148226
rect 497214 148170 497282 148226
rect 497338 148170 497406 148226
rect 497462 148170 497558 148226
rect 496938 148102 497558 148170
rect 496938 148046 497034 148102
rect 497090 148046 497158 148102
rect 497214 148046 497282 148102
rect 497338 148046 497406 148102
rect 497462 148046 497558 148102
rect 496938 147978 497558 148046
rect 496938 147922 497034 147978
rect 497090 147922 497158 147978
rect 497214 147922 497282 147978
rect 497338 147922 497406 147978
rect 497462 147922 497558 147978
rect 471996 142318 472052 142328
rect 471996 141988 472052 142262
rect 471996 141922 472052 141932
rect 484428 141958 484484 141968
rect 484428 141764 484484 141902
rect 484428 141698 484484 141708
rect 469938 136294 470034 136350
rect 470090 136294 470158 136350
rect 470214 136294 470282 136350
rect 470338 136294 470406 136350
rect 470462 136294 470558 136350
rect 469938 136226 470558 136294
rect 469938 136170 470034 136226
rect 470090 136170 470158 136226
rect 470214 136170 470282 136226
rect 470338 136170 470406 136226
rect 470462 136170 470558 136226
rect 469938 136102 470558 136170
rect 469938 136046 470034 136102
rect 470090 136046 470158 136102
rect 470214 136046 470282 136102
rect 470338 136046 470406 136102
rect 470462 136046 470558 136102
rect 469938 135978 470558 136046
rect 469938 135922 470034 135978
rect 470090 135922 470158 135978
rect 470214 135922 470282 135978
rect 470338 135922 470406 135978
rect 470462 135922 470558 135978
rect 469938 118350 470558 135922
rect 469938 118294 470034 118350
rect 470090 118294 470158 118350
rect 470214 118294 470282 118350
rect 470338 118294 470406 118350
rect 470462 118294 470558 118350
rect 469938 118226 470558 118294
rect 469938 118170 470034 118226
rect 470090 118170 470158 118226
rect 470214 118170 470282 118226
rect 470338 118170 470406 118226
rect 470462 118170 470558 118226
rect 469938 118102 470558 118170
rect 469938 118046 470034 118102
rect 470090 118046 470158 118102
rect 470214 118046 470282 118102
rect 470338 118046 470406 118102
rect 470462 118046 470558 118102
rect 469938 117978 470558 118046
rect 469938 117922 470034 117978
rect 470090 117922 470158 117978
rect 470214 117922 470282 117978
rect 470338 117922 470406 117978
rect 470462 117922 470558 117978
rect 469938 100350 470558 117922
rect 469938 100294 470034 100350
rect 470090 100294 470158 100350
rect 470214 100294 470282 100350
rect 470338 100294 470406 100350
rect 470462 100294 470558 100350
rect 469938 100226 470558 100294
rect 469938 100170 470034 100226
rect 470090 100170 470158 100226
rect 470214 100170 470282 100226
rect 470338 100170 470406 100226
rect 470462 100170 470558 100226
rect 469938 100102 470558 100170
rect 469938 100046 470034 100102
rect 470090 100046 470158 100102
rect 470214 100046 470282 100102
rect 470338 100046 470406 100102
rect 470462 100046 470558 100102
rect 469938 99978 470558 100046
rect 469938 99922 470034 99978
rect 470090 99922 470158 99978
rect 470214 99922 470282 99978
rect 470338 99922 470406 99978
rect 470462 99922 470558 99978
rect 469938 82350 470558 99922
rect 469938 82294 470034 82350
rect 470090 82294 470158 82350
rect 470214 82294 470282 82350
rect 470338 82294 470406 82350
rect 470462 82294 470558 82350
rect 469938 82226 470558 82294
rect 469938 82170 470034 82226
rect 470090 82170 470158 82226
rect 470214 82170 470282 82226
rect 470338 82170 470406 82226
rect 470462 82170 470558 82226
rect 469938 82102 470558 82170
rect 469938 82046 470034 82102
rect 470090 82046 470158 82102
rect 470214 82046 470282 82102
rect 470338 82046 470406 82102
rect 470462 82046 470558 82102
rect 469938 81978 470558 82046
rect 469938 81922 470034 81978
rect 470090 81922 470158 81978
rect 470214 81922 470282 81978
rect 470338 81922 470406 81978
rect 470462 81922 470558 81978
rect 469938 64350 470558 81922
rect 469938 64294 470034 64350
rect 470090 64294 470158 64350
rect 470214 64294 470282 64350
rect 470338 64294 470406 64350
rect 470462 64294 470558 64350
rect 469938 64226 470558 64294
rect 469938 64170 470034 64226
rect 470090 64170 470158 64226
rect 470214 64170 470282 64226
rect 470338 64170 470406 64226
rect 470462 64170 470558 64226
rect 469938 64102 470558 64170
rect 469938 64046 470034 64102
rect 470090 64046 470158 64102
rect 470214 64046 470282 64102
rect 470338 64046 470406 64102
rect 470462 64046 470558 64102
rect 469938 63978 470558 64046
rect 469938 63922 470034 63978
rect 470090 63922 470158 63978
rect 470214 63922 470282 63978
rect 470338 63922 470406 63978
rect 470462 63922 470558 63978
rect 469938 46350 470558 63922
rect 469938 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 470558 46350
rect 469938 46226 470558 46294
rect 469938 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 470558 46226
rect 469938 46102 470558 46170
rect 469938 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 470558 46102
rect 469938 45978 470558 46046
rect 469938 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 470558 45978
rect 469938 28350 470558 45922
rect 469938 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 470558 28350
rect 469938 28226 470558 28294
rect 469938 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 470558 28226
rect 469938 28102 470558 28170
rect 469938 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 470558 28102
rect 469938 27978 470558 28046
rect 469938 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 470558 27978
rect 469938 10350 470558 27922
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 469938 -1120 470558 9922
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 130350 497558 147922
rect 500658 298350 501278 305970
rect 500658 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 501278 298350
rect 500658 298226 501278 298294
rect 500658 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 501278 298226
rect 500658 298102 501278 298170
rect 500658 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 501278 298102
rect 500658 297978 501278 298046
rect 500658 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 501278 297978
rect 500658 280350 501278 297922
rect 500658 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 501278 280350
rect 500658 280226 501278 280294
rect 500658 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 501278 280226
rect 500658 280102 501278 280170
rect 500658 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 501278 280102
rect 500658 279978 501278 280046
rect 500658 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 501278 279978
rect 500658 262350 501278 279922
rect 500658 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 501278 262350
rect 500658 262226 501278 262294
rect 500658 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 501278 262226
rect 500658 262102 501278 262170
rect 500658 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 501278 262102
rect 500658 261978 501278 262046
rect 500658 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 501278 261978
rect 500658 244350 501278 261922
rect 500658 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 501278 244350
rect 500658 244226 501278 244294
rect 500658 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 501278 244226
rect 500658 244102 501278 244170
rect 500658 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 501278 244102
rect 500658 243978 501278 244046
rect 500658 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 501278 243978
rect 500658 226350 501278 243922
rect 500658 226294 500754 226350
rect 500810 226294 500878 226350
rect 500934 226294 501002 226350
rect 501058 226294 501126 226350
rect 501182 226294 501278 226350
rect 500658 226226 501278 226294
rect 500658 226170 500754 226226
rect 500810 226170 500878 226226
rect 500934 226170 501002 226226
rect 501058 226170 501126 226226
rect 501182 226170 501278 226226
rect 500658 226102 501278 226170
rect 500658 226046 500754 226102
rect 500810 226046 500878 226102
rect 500934 226046 501002 226102
rect 501058 226046 501126 226102
rect 501182 226046 501278 226102
rect 500658 225978 501278 226046
rect 500658 225922 500754 225978
rect 500810 225922 500878 225978
rect 500934 225922 501002 225978
rect 501058 225922 501126 225978
rect 501182 225922 501278 225978
rect 500658 208350 501278 225922
rect 500658 208294 500754 208350
rect 500810 208294 500878 208350
rect 500934 208294 501002 208350
rect 501058 208294 501126 208350
rect 501182 208294 501278 208350
rect 500658 208226 501278 208294
rect 500658 208170 500754 208226
rect 500810 208170 500878 208226
rect 500934 208170 501002 208226
rect 501058 208170 501126 208226
rect 501182 208170 501278 208226
rect 500658 208102 501278 208170
rect 500658 208046 500754 208102
rect 500810 208046 500878 208102
rect 500934 208046 501002 208102
rect 501058 208046 501126 208102
rect 501182 208046 501278 208102
rect 500658 207978 501278 208046
rect 500658 207922 500754 207978
rect 500810 207922 500878 207978
rect 500934 207922 501002 207978
rect 501058 207922 501126 207978
rect 501182 207922 501278 207978
rect 500658 190350 501278 207922
rect 500658 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 501278 190350
rect 500658 190226 501278 190294
rect 500658 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 501278 190226
rect 500658 190102 501278 190170
rect 500658 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 501278 190102
rect 500658 189978 501278 190046
rect 500658 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 501278 189978
rect 500658 172350 501278 189922
rect 500658 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 501278 172350
rect 500658 172226 501278 172294
rect 500658 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 501278 172226
rect 500658 172102 501278 172170
rect 500658 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 501278 172102
rect 500658 171978 501278 172046
rect 500658 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 501278 171978
rect 500658 154350 501278 171922
rect 500658 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 501278 154350
rect 500658 154226 501278 154294
rect 500658 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 501278 154226
rect 500658 154102 501278 154170
rect 500658 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 501278 154102
rect 500658 153978 501278 154046
rect 500658 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 501278 153978
rect 498988 142884 499044 142894
rect 498988 142678 499044 142828
rect 498988 142612 499044 142622
rect 496938 130294 497034 130350
rect 497090 130294 497158 130350
rect 497214 130294 497282 130350
rect 497338 130294 497406 130350
rect 497462 130294 497558 130350
rect 496938 130226 497558 130294
rect 496938 130170 497034 130226
rect 497090 130170 497158 130226
rect 497214 130170 497282 130226
rect 497338 130170 497406 130226
rect 497462 130170 497558 130226
rect 496938 130102 497558 130170
rect 496938 130046 497034 130102
rect 497090 130046 497158 130102
rect 497214 130046 497282 130102
rect 497338 130046 497406 130102
rect 497462 130046 497558 130102
rect 496938 129978 497558 130046
rect 496938 129922 497034 129978
rect 497090 129922 497158 129978
rect 497214 129922 497282 129978
rect 497338 129922 497406 129978
rect 497462 129922 497558 129978
rect 496938 112350 497558 129922
rect 496938 112294 497034 112350
rect 497090 112294 497158 112350
rect 497214 112294 497282 112350
rect 497338 112294 497406 112350
rect 497462 112294 497558 112350
rect 496938 112226 497558 112294
rect 496938 112170 497034 112226
rect 497090 112170 497158 112226
rect 497214 112170 497282 112226
rect 497338 112170 497406 112226
rect 497462 112170 497558 112226
rect 496938 112102 497558 112170
rect 496938 112046 497034 112102
rect 497090 112046 497158 112102
rect 497214 112046 497282 112102
rect 497338 112046 497406 112102
rect 497462 112046 497558 112102
rect 496938 111978 497558 112046
rect 496938 111922 497034 111978
rect 497090 111922 497158 111978
rect 497214 111922 497282 111978
rect 497338 111922 497406 111978
rect 497462 111922 497558 111978
rect 496938 94350 497558 111922
rect 496938 94294 497034 94350
rect 497090 94294 497158 94350
rect 497214 94294 497282 94350
rect 497338 94294 497406 94350
rect 497462 94294 497558 94350
rect 496938 94226 497558 94294
rect 496938 94170 497034 94226
rect 497090 94170 497158 94226
rect 497214 94170 497282 94226
rect 497338 94170 497406 94226
rect 497462 94170 497558 94226
rect 496938 94102 497558 94170
rect 496938 94046 497034 94102
rect 497090 94046 497158 94102
rect 497214 94046 497282 94102
rect 497338 94046 497406 94102
rect 497462 94046 497558 94102
rect 496938 93978 497558 94046
rect 496938 93922 497034 93978
rect 497090 93922 497158 93978
rect 497214 93922 497282 93978
rect 497338 93922 497406 93978
rect 497462 93922 497558 93978
rect 496938 76350 497558 93922
rect 496938 76294 497034 76350
rect 497090 76294 497158 76350
rect 497214 76294 497282 76350
rect 497338 76294 497406 76350
rect 497462 76294 497558 76350
rect 496938 76226 497558 76294
rect 496938 76170 497034 76226
rect 497090 76170 497158 76226
rect 497214 76170 497282 76226
rect 497338 76170 497406 76226
rect 497462 76170 497558 76226
rect 496938 76102 497558 76170
rect 496938 76046 497034 76102
rect 497090 76046 497158 76102
rect 497214 76046 497282 76102
rect 497338 76046 497406 76102
rect 497462 76046 497558 76102
rect 496938 75978 497558 76046
rect 496938 75922 497034 75978
rect 497090 75922 497158 75978
rect 497214 75922 497282 75978
rect 497338 75922 497406 75978
rect 497462 75922 497558 75978
rect 496938 58350 497558 75922
rect 496938 58294 497034 58350
rect 497090 58294 497158 58350
rect 497214 58294 497282 58350
rect 497338 58294 497406 58350
rect 497462 58294 497558 58350
rect 496938 58226 497558 58294
rect 496938 58170 497034 58226
rect 497090 58170 497158 58226
rect 497214 58170 497282 58226
rect 497338 58170 497406 58226
rect 497462 58170 497558 58226
rect 496938 58102 497558 58170
rect 496938 58046 497034 58102
rect 497090 58046 497158 58102
rect 497214 58046 497282 58102
rect 497338 58046 497406 58102
rect 497462 58046 497558 58102
rect 496938 57978 497558 58046
rect 496938 57922 497034 57978
rect 497090 57922 497158 57978
rect 497214 57922 497282 57978
rect 497338 57922 497406 57978
rect 497462 57922 497558 57978
rect 496938 40350 497558 57922
rect 496938 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 497558 40350
rect 496938 40226 497558 40294
rect 496938 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 497558 40226
rect 496938 40102 497558 40170
rect 496938 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 497558 40102
rect 496938 39978 497558 40046
rect 496938 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 497558 39978
rect 496938 22350 497558 39922
rect 496938 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 497558 22350
rect 496938 22226 497558 22294
rect 496938 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 497558 22226
rect 496938 22102 497558 22170
rect 496938 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 497558 22102
rect 496938 21978 497558 22046
rect 496938 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 497558 21978
rect 496938 4350 497558 21922
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 496938 -160 497558 3922
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 136350 501278 153922
rect 527658 292350 528278 309922
rect 527658 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 528278 292350
rect 527658 292226 528278 292294
rect 527658 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 528278 292226
rect 527658 292102 528278 292170
rect 527658 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 528278 292102
rect 527658 291978 528278 292046
rect 527658 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 528278 291978
rect 527658 274350 528278 291922
rect 527658 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 528278 274350
rect 527658 274226 528278 274294
rect 527658 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 528278 274226
rect 527658 274102 528278 274170
rect 527658 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 528278 274102
rect 527658 273978 528278 274046
rect 527658 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 528278 273978
rect 527658 256350 528278 273922
rect 527658 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 528278 256350
rect 527658 256226 528278 256294
rect 527658 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 528278 256226
rect 527658 256102 528278 256170
rect 527658 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 528278 256102
rect 527658 255978 528278 256046
rect 527658 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255922 528278 255978
rect 527658 238350 528278 255922
rect 527658 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 528278 238350
rect 527658 238226 528278 238294
rect 527658 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 528278 238226
rect 527658 238102 528278 238170
rect 527658 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 528278 238102
rect 527658 237978 528278 238046
rect 527658 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 528278 237978
rect 527658 220350 528278 237922
rect 527658 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 528278 220350
rect 527658 220226 528278 220294
rect 527658 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 528278 220226
rect 527658 220102 528278 220170
rect 527658 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 528278 220102
rect 527658 219978 528278 220046
rect 527658 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 528278 219978
rect 527658 202350 528278 219922
rect 527658 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 528278 202350
rect 527658 202226 528278 202294
rect 527658 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 528278 202226
rect 527658 202102 528278 202170
rect 527658 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 528278 202102
rect 527658 201978 528278 202046
rect 527658 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 528278 201978
rect 527658 184350 528278 201922
rect 527658 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 528278 184350
rect 527658 184226 528278 184294
rect 527658 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 528278 184226
rect 527658 184102 528278 184170
rect 527658 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 528278 184102
rect 527658 183978 528278 184046
rect 527658 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 528278 183978
rect 527658 166350 528278 183922
rect 527658 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 528278 166350
rect 527658 166226 528278 166294
rect 527658 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 528278 166226
rect 527658 166102 528278 166170
rect 527658 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 528278 166102
rect 527658 165978 528278 166046
rect 527658 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 528278 165978
rect 527658 148350 528278 165922
rect 527658 148294 527754 148350
rect 527810 148294 527878 148350
rect 527934 148294 528002 148350
rect 528058 148294 528126 148350
rect 528182 148294 528278 148350
rect 527658 148226 528278 148294
rect 527658 148170 527754 148226
rect 527810 148170 527878 148226
rect 527934 148170 528002 148226
rect 528058 148170 528126 148226
rect 528182 148170 528278 148226
rect 527658 148102 528278 148170
rect 527658 148046 527754 148102
rect 527810 148046 527878 148102
rect 527934 148046 528002 148102
rect 528058 148046 528126 148102
rect 528182 148046 528278 148102
rect 527658 147978 528278 148046
rect 527658 147922 527754 147978
rect 527810 147922 527878 147978
rect 527934 147922 528002 147978
rect 528058 147922 528126 147978
rect 528182 147922 528278 147978
rect 505596 141540 505652 141550
rect 505596 141058 505652 141484
rect 505596 140992 505652 141002
rect 500658 136294 500754 136350
rect 500810 136294 500878 136350
rect 500934 136294 501002 136350
rect 501058 136294 501126 136350
rect 501182 136294 501278 136350
rect 500658 136226 501278 136294
rect 500658 136170 500754 136226
rect 500810 136170 500878 136226
rect 500934 136170 501002 136226
rect 501058 136170 501126 136226
rect 501182 136170 501278 136226
rect 500658 136102 501278 136170
rect 500658 136046 500754 136102
rect 500810 136046 500878 136102
rect 500934 136046 501002 136102
rect 501058 136046 501126 136102
rect 501182 136046 501278 136102
rect 500658 135978 501278 136046
rect 500658 135922 500754 135978
rect 500810 135922 500878 135978
rect 500934 135922 501002 135978
rect 501058 135922 501126 135978
rect 501182 135922 501278 135978
rect 500658 118350 501278 135922
rect 500658 118294 500754 118350
rect 500810 118294 500878 118350
rect 500934 118294 501002 118350
rect 501058 118294 501126 118350
rect 501182 118294 501278 118350
rect 500658 118226 501278 118294
rect 500658 118170 500754 118226
rect 500810 118170 500878 118226
rect 500934 118170 501002 118226
rect 501058 118170 501126 118226
rect 501182 118170 501278 118226
rect 500658 118102 501278 118170
rect 500658 118046 500754 118102
rect 500810 118046 500878 118102
rect 500934 118046 501002 118102
rect 501058 118046 501126 118102
rect 501182 118046 501278 118102
rect 500658 117978 501278 118046
rect 500658 117922 500754 117978
rect 500810 117922 500878 117978
rect 500934 117922 501002 117978
rect 501058 117922 501126 117978
rect 501182 117922 501278 117978
rect 500658 100350 501278 117922
rect 500658 100294 500754 100350
rect 500810 100294 500878 100350
rect 500934 100294 501002 100350
rect 501058 100294 501126 100350
rect 501182 100294 501278 100350
rect 500658 100226 501278 100294
rect 500658 100170 500754 100226
rect 500810 100170 500878 100226
rect 500934 100170 501002 100226
rect 501058 100170 501126 100226
rect 501182 100170 501278 100226
rect 500658 100102 501278 100170
rect 500658 100046 500754 100102
rect 500810 100046 500878 100102
rect 500934 100046 501002 100102
rect 501058 100046 501126 100102
rect 501182 100046 501278 100102
rect 500658 99978 501278 100046
rect 500658 99922 500754 99978
rect 500810 99922 500878 99978
rect 500934 99922 501002 99978
rect 501058 99922 501126 99978
rect 501182 99922 501278 99978
rect 500658 82350 501278 99922
rect 500658 82294 500754 82350
rect 500810 82294 500878 82350
rect 500934 82294 501002 82350
rect 501058 82294 501126 82350
rect 501182 82294 501278 82350
rect 500658 82226 501278 82294
rect 500658 82170 500754 82226
rect 500810 82170 500878 82226
rect 500934 82170 501002 82226
rect 501058 82170 501126 82226
rect 501182 82170 501278 82226
rect 500658 82102 501278 82170
rect 500658 82046 500754 82102
rect 500810 82046 500878 82102
rect 500934 82046 501002 82102
rect 501058 82046 501126 82102
rect 501182 82046 501278 82102
rect 500658 81978 501278 82046
rect 500658 81922 500754 81978
rect 500810 81922 500878 81978
rect 500934 81922 501002 81978
rect 501058 81922 501126 81978
rect 501182 81922 501278 81978
rect 500658 64350 501278 81922
rect 500658 64294 500754 64350
rect 500810 64294 500878 64350
rect 500934 64294 501002 64350
rect 501058 64294 501126 64350
rect 501182 64294 501278 64350
rect 500658 64226 501278 64294
rect 500658 64170 500754 64226
rect 500810 64170 500878 64226
rect 500934 64170 501002 64226
rect 501058 64170 501126 64226
rect 501182 64170 501278 64226
rect 500658 64102 501278 64170
rect 500658 64046 500754 64102
rect 500810 64046 500878 64102
rect 500934 64046 501002 64102
rect 501058 64046 501126 64102
rect 501182 64046 501278 64102
rect 500658 63978 501278 64046
rect 500658 63922 500754 63978
rect 500810 63922 500878 63978
rect 500934 63922 501002 63978
rect 501058 63922 501126 63978
rect 501182 63922 501278 63978
rect 500658 46350 501278 63922
rect 500658 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 501278 46350
rect 500658 46226 501278 46294
rect 500658 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 501278 46226
rect 500658 46102 501278 46170
rect 500658 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 501278 46102
rect 500658 45978 501278 46046
rect 500658 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 501278 45978
rect 500658 28350 501278 45922
rect 500658 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 501278 28350
rect 500658 28226 501278 28294
rect 500658 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 501278 28226
rect 500658 28102 501278 28170
rect 500658 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 501278 28102
rect 500658 27978 501278 28046
rect 500658 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 501278 27978
rect 500658 10350 501278 27922
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 500658 -1120 501278 9922
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 130350 528278 147922
rect 527658 130294 527754 130350
rect 527810 130294 527878 130350
rect 527934 130294 528002 130350
rect 528058 130294 528126 130350
rect 528182 130294 528278 130350
rect 527658 130226 528278 130294
rect 527658 130170 527754 130226
rect 527810 130170 527878 130226
rect 527934 130170 528002 130226
rect 528058 130170 528126 130226
rect 528182 130170 528278 130226
rect 527658 130102 528278 130170
rect 527658 130046 527754 130102
rect 527810 130046 527878 130102
rect 527934 130046 528002 130102
rect 528058 130046 528126 130102
rect 528182 130046 528278 130102
rect 527658 129978 528278 130046
rect 527658 129922 527754 129978
rect 527810 129922 527878 129978
rect 527934 129922 528002 129978
rect 528058 129922 528126 129978
rect 528182 129922 528278 129978
rect 527658 112350 528278 129922
rect 527658 112294 527754 112350
rect 527810 112294 527878 112350
rect 527934 112294 528002 112350
rect 528058 112294 528126 112350
rect 528182 112294 528278 112350
rect 527658 112226 528278 112294
rect 527658 112170 527754 112226
rect 527810 112170 527878 112226
rect 527934 112170 528002 112226
rect 528058 112170 528126 112226
rect 528182 112170 528278 112226
rect 527658 112102 528278 112170
rect 527658 112046 527754 112102
rect 527810 112046 527878 112102
rect 527934 112046 528002 112102
rect 528058 112046 528126 112102
rect 528182 112046 528278 112102
rect 527658 111978 528278 112046
rect 527658 111922 527754 111978
rect 527810 111922 527878 111978
rect 527934 111922 528002 111978
rect 528058 111922 528126 111978
rect 528182 111922 528278 111978
rect 527658 94350 528278 111922
rect 527658 94294 527754 94350
rect 527810 94294 527878 94350
rect 527934 94294 528002 94350
rect 528058 94294 528126 94350
rect 528182 94294 528278 94350
rect 527658 94226 528278 94294
rect 527658 94170 527754 94226
rect 527810 94170 527878 94226
rect 527934 94170 528002 94226
rect 528058 94170 528126 94226
rect 528182 94170 528278 94226
rect 527658 94102 528278 94170
rect 527658 94046 527754 94102
rect 527810 94046 527878 94102
rect 527934 94046 528002 94102
rect 528058 94046 528126 94102
rect 528182 94046 528278 94102
rect 527658 93978 528278 94046
rect 527658 93922 527754 93978
rect 527810 93922 527878 93978
rect 527934 93922 528002 93978
rect 528058 93922 528126 93978
rect 528182 93922 528278 93978
rect 527658 76350 528278 93922
rect 527658 76294 527754 76350
rect 527810 76294 527878 76350
rect 527934 76294 528002 76350
rect 528058 76294 528126 76350
rect 528182 76294 528278 76350
rect 527658 76226 528278 76294
rect 527658 76170 527754 76226
rect 527810 76170 527878 76226
rect 527934 76170 528002 76226
rect 528058 76170 528126 76226
rect 528182 76170 528278 76226
rect 527658 76102 528278 76170
rect 527658 76046 527754 76102
rect 527810 76046 527878 76102
rect 527934 76046 528002 76102
rect 528058 76046 528126 76102
rect 528182 76046 528278 76102
rect 527658 75978 528278 76046
rect 527658 75922 527754 75978
rect 527810 75922 527878 75978
rect 527934 75922 528002 75978
rect 528058 75922 528126 75978
rect 528182 75922 528278 75978
rect 527658 58350 528278 75922
rect 527658 58294 527754 58350
rect 527810 58294 527878 58350
rect 527934 58294 528002 58350
rect 528058 58294 528126 58350
rect 528182 58294 528278 58350
rect 527658 58226 528278 58294
rect 527658 58170 527754 58226
rect 527810 58170 527878 58226
rect 527934 58170 528002 58226
rect 528058 58170 528126 58226
rect 528182 58170 528278 58226
rect 527658 58102 528278 58170
rect 527658 58046 527754 58102
rect 527810 58046 527878 58102
rect 527934 58046 528002 58102
rect 528058 58046 528126 58102
rect 528182 58046 528278 58102
rect 527658 57978 528278 58046
rect 527658 57922 527754 57978
rect 527810 57922 527878 57978
rect 527934 57922 528002 57978
rect 528058 57922 528126 57978
rect 528182 57922 528278 57978
rect 527658 40350 528278 57922
rect 527658 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 528278 40350
rect 527658 40226 528278 40294
rect 527658 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 528278 40226
rect 527658 40102 528278 40170
rect 527658 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 528278 40102
rect 527658 39978 528278 40046
rect 527658 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 528278 39978
rect 527658 22350 528278 39922
rect 527658 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 528278 22350
rect 527658 22226 528278 22294
rect 527658 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 528278 22226
rect 527658 22102 528278 22170
rect 527658 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 528278 22102
rect 527658 21978 528278 22046
rect 527658 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 528278 21978
rect 527658 4350 528278 21922
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 442350 531998 453058
rect 533036 451556 533092 451566
rect 533036 450212 533092 451500
rect 533036 450146 533092 450156
rect 531378 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 531998 442350
rect 531378 442226 531998 442294
rect 531378 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 531998 442226
rect 531378 442102 531998 442170
rect 531378 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 531998 442102
rect 531378 441978 531998 442046
rect 531378 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 531998 441978
rect 531378 424350 531998 441922
rect 531378 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 531998 424350
rect 531378 424226 531998 424294
rect 531378 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 531998 424226
rect 531378 424102 531998 424170
rect 531378 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 531998 424102
rect 531378 423978 531998 424046
rect 531378 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 531998 423978
rect 531378 406350 531998 423922
rect 531378 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 531998 406350
rect 531378 406226 531998 406294
rect 531378 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 531998 406226
rect 531378 406102 531998 406170
rect 531378 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 531998 406102
rect 531378 405978 531998 406046
rect 531378 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 531998 405978
rect 531378 388350 531998 405922
rect 548156 390628 548212 537740
rect 549388 536004 549444 536014
rect 549388 394212 549444 535948
rect 549500 533428 549556 533438
rect 549500 399588 549556 533372
rect 556108 518868 556164 546182
rect 556220 529396 556276 546362
rect 556220 529330 556276 529340
rect 558378 544350 558998 561922
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 556108 518802 556164 518812
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 551248 514350 551568 514384
rect 551248 514294 551318 514350
rect 551374 514294 551442 514350
rect 551498 514294 551568 514350
rect 551248 514226 551568 514294
rect 551248 514170 551318 514226
rect 551374 514170 551442 514226
rect 551498 514170 551568 514226
rect 551248 514102 551568 514170
rect 551248 514046 551318 514102
rect 551374 514046 551442 514102
rect 551498 514046 551568 514102
rect 551248 513978 551568 514046
rect 551248 513922 551318 513978
rect 551374 513922 551442 513978
rect 551498 513922 551568 513978
rect 551248 513888 551568 513922
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 551248 496350 551568 496384
rect 551248 496294 551318 496350
rect 551374 496294 551442 496350
rect 551498 496294 551568 496350
rect 551248 496226 551568 496294
rect 551248 496170 551318 496226
rect 551374 496170 551442 496226
rect 551498 496170 551568 496226
rect 551248 496102 551568 496170
rect 551248 496046 551318 496102
rect 551374 496046 551442 496102
rect 551498 496046 551568 496102
rect 551248 495978 551568 496046
rect 551248 495922 551318 495978
rect 551374 495922 551442 495978
rect 551498 495922 551568 495978
rect 551248 495888 551568 495922
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 551248 478350 551568 478384
rect 551248 478294 551318 478350
rect 551374 478294 551442 478350
rect 551498 478294 551568 478350
rect 551248 478226 551568 478294
rect 551248 478170 551318 478226
rect 551374 478170 551442 478226
rect 551498 478170 551568 478226
rect 551248 478102 551568 478170
rect 551248 478046 551318 478102
rect 551374 478046 551442 478102
rect 551498 478046 551568 478102
rect 551248 477978 551568 478046
rect 551248 477922 551318 477978
rect 551374 477922 551442 477978
rect 551498 477922 551568 477978
rect 551248 477888 551568 477922
rect 558378 472350 558998 489922
rect 558378 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 558998 472350
rect 558378 472226 558998 472294
rect 558378 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 558998 472226
rect 558378 472102 558998 472170
rect 558378 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 558998 472102
rect 558378 471978 558998 472046
rect 558378 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 558998 471978
rect 551248 460350 551568 460384
rect 551248 460294 551318 460350
rect 551374 460294 551442 460350
rect 551498 460294 551568 460350
rect 551248 460226 551568 460294
rect 551248 460170 551318 460226
rect 551374 460170 551442 460226
rect 551498 460170 551568 460226
rect 551248 460102 551568 460170
rect 551248 460046 551318 460102
rect 551374 460046 551442 460102
rect 551498 460046 551568 460102
rect 551248 459978 551568 460046
rect 551248 459922 551318 459978
rect 551374 459922 551442 459978
rect 551498 459922 551568 459978
rect 551248 459888 551568 459922
rect 554428 455252 554484 455262
rect 554428 450436 554484 455196
rect 554428 450370 554484 450380
rect 558378 454350 558998 471922
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 549500 399522 549556 399532
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 558378 400350 558998 417922
rect 558378 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 558998 400350
rect 558378 400226 558998 400294
rect 558378 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 558998 400226
rect 558378 400102 558998 400170
rect 558378 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 558998 400102
rect 558378 399978 558998 400046
rect 558378 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 558998 399978
rect 549388 394146 549444 394156
rect 548156 390562 548212 390572
rect 531378 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388294 531998 388350
rect 531378 388226 531998 388294
rect 531378 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 531998 388226
rect 531378 388102 531998 388170
rect 531378 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 531998 388102
rect 531378 387978 531998 388046
rect 531378 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 531998 387978
rect 531378 370350 531998 387922
rect 531378 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 531998 370350
rect 531378 370226 531998 370294
rect 531378 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 531998 370226
rect 531378 370102 531998 370170
rect 531378 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 531998 370102
rect 531378 369978 531998 370046
rect 531378 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 531998 369978
rect 531378 352350 531998 369922
rect 531378 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 531998 352350
rect 531378 352226 531998 352294
rect 531378 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 531998 352226
rect 531378 352102 531998 352170
rect 531378 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 531998 352102
rect 531378 351978 531998 352046
rect 531378 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 531998 351978
rect 531378 334350 531998 351922
rect 531378 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 531998 334350
rect 531378 334226 531998 334294
rect 531378 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 531998 334226
rect 531378 334102 531998 334170
rect 531378 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 531998 334102
rect 531378 333978 531998 334046
rect 531378 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 531998 333978
rect 531378 316350 531998 333922
rect 531378 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 531998 316350
rect 531378 316226 531998 316294
rect 531378 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 531998 316226
rect 531378 316102 531998 316170
rect 531378 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 531998 316102
rect 531378 315978 531998 316046
rect 531378 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 531998 315978
rect 531378 298350 531998 315922
rect 531378 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 531998 298350
rect 531378 298226 531998 298294
rect 531378 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 531998 298226
rect 531378 298102 531998 298170
rect 531378 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 531998 298102
rect 531378 297978 531998 298046
rect 531378 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 531998 297978
rect 531378 280350 531998 297922
rect 531378 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 531998 280350
rect 531378 280226 531998 280294
rect 531378 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 531998 280226
rect 531378 280102 531998 280170
rect 531378 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 531998 280102
rect 531378 279978 531998 280046
rect 531378 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 531998 279978
rect 531378 262350 531998 279922
rect 531378 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 531998 262350
rect 531378 262226 531998 262294
rect 531378 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 531998 262226
rect 531378 262102 531998 262170
rect 531378 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 531998 262102
rect 531378 261978 531998 262046
rect 531378 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 531998 261978
rect 531378 244350 531998 261922
rect 558378 382350 558998 399922
rect 558378 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 558998 382350
rect 558378 382226 558998 382294
rect 558378 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 558998 382226
rect 558378 382102 558998 382170
rect 558378 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 558998 382102
rect 558378 381978 558998 382046
rect 558378 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 558998 381978
rect 558378 364350 558998 381922
rect 558378 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 558998 364350
rect 558378 364226 558998 364294
rect 558378 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 558998 364226
rect 558378 364102 558998 364170
rect 558378 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 558998 364102
rect 558378 363978 558998 364046
rect 558378 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 558998 363978
rect 558378 346350 558998 363922
rect 558378 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 558998 346350
rect 558378 346226 558998 346294
rect 558378 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 558998 346226
rect 558378 346102 558998 346170
rect 558378 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 558998 346102
rect 558378 345978 558998 346046
rect 558378 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 558998 345978
rect 558378 328350 558998 345922
rect 558378 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 558998 328350
rect 558378 328226 558998 328294
rect 558378 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 558998 328226
rect 558378 328102 558998 328170
rect 558378 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 558998 328102
rect 558378 327978 558998 328046
rect 558378 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 558998 327978
rect 558378 310350 558998 327922
rect 558378 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 558998 310350
rect 558378 310226 558998 310294
rect 558378 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 558998 310226
rect 558378 310102 558998 310170
rect 558378 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 558998 310102
rect 558378 309978 558998 310046
rect 558378 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 558998 309978
rect 558378 292350 558998 309922
rect 558378 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 558998 292350
rect 558378 292226 558998 292294
rect 558378 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 558998 292226
rect 558378 292102 558998 292170
rect 558378 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 558998 292102
rect 558378 291978 558998 292046
rect 558378 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 558998 291978
rect 558378 274350 558998 291922
rect 558378 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 558998 274350
rect 558378 274226 558998 274294
rect 558378 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 558998 274226
rect 558378 274102 558998 274170
rect 558378 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 558998 274102
rect 558378 273978 558998 274046
rect 558378 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 558998 273978
rect 558378 256350 558998 273922
rect 558378 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 558998 256350
rect 558378 256226 558998 256294
rect 558378 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 558998 256226
rect 558378 256102 558998 256170
rect 558378 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 558998 256102
rect 557390 256023 557866 256040
rect 557390 255967 557414 256023
rect 557470 255967 557538 256023
rect 557594 255967 557662 256023
rect 557718 255967 557786 256023
rect 557842 255967 557866 256023
rect 557390 255899 557866 255967
rect 557390 255843 557414 255899
rect 557470 255843 557538 255899
rect 557594 255843 557662 255899
rect 557718 255843 557786 255899
rect 557842 255843 557866 255899
rect 557390 255826 557866 255843
rect 558378 255978 558998 256046
rect 558378 255922 558474 255978
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 558998 255978
rect 531378 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 531998 244350
rect 531378 244226 531998 244294
rect 531378 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 531998 244226
rect 531378 244102 531998 244170
rect 531378 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 531998 244102
rect 531378 243978 531998 244046
rect 531378 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 531998 243978
rect 531378 226350 531998 243922
rect 556590 244350 557066 244384
rect 556590 244294 556614 244350
rect 556670 244294 556738 244350
rect 556794 244294 556862 244350
rect 556918 244294 556986 244350
rect 557042 244294 557066 244350
rect 556590 244226 557066 244294
rect 556590 244170 556614 244226
rect 556670 244170 556738 244226
rect 556794 244170 556862 244226
rect 556918 244170 556986 244226
rect 557042 244170 557066 244226
rect 556590 244102 557066 244170
rect 556590 244046 556614 244102
rect 556670 244046 556738 244102
rect 556794 244046 556862 244102
rect 556918 244046 556986 244102
rect 557042 244046 557066 244102
rect 556590 243978 557066 244046
rect 556590 243922 556614 243978
rect 556670 243922 556738 243978
rect 556794 243922 556862 243978
rect 556918 243922 556986 243978
rect 557042 243922 557066 243978
rect 556590 243888 557066 243922
rect 557390 238350 557866 238384
rect 557390 238294 557414 238350
rect 557470 238294 557538 238350
rect 557594 238294 557662 238350
rect 557718 238294 557786 238350
rect 557842 238294 557866 238350
rect 557390 238226 557866 238294
rect 557390 238170 557414 238226
rect 557470 238170 557538 238226
rect 557594 238170 557662 238226
rect 557718 238170 557786 238226
rect 557842 238170 557866 238226
rect 557390 238102 557866 238170
rect 557390 238046 557414 238102
rect 557470 238046 557538 238102
rect 557594 238046 557662 238102
rect 557718 238046 557786 238102
rect 557842 238046 557866 238102
rect 557390 237978 557866 238046
rect 557390 237922 557414 237978
rect 557470 237922 557538 237978
rect 557594 237922 557662 237978
rect 557718 237922 557786 237978
rect 557842 237922 557866 237978
rect 557390 237888 557866 237922
rect 558378 238350 558998 255922
rect 558378 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 558998 238350
rect 558378 238226 558998 238294
rect 558378 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 558998 238226
rect 558378 238102 558998 238170
rect 558378 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 558998 238102
rect 558378 237978 558998 238046
rect 558378 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 558998 237978
rect 531378 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 531998 226350
rect 531378 226226 531998 226294
rect 531378 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 531998 226226
rect 531378 226102 531998 226170
rect 531378 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 531998 226102
rect 531378 225978 531998 226046
rect 531378 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 531998 225978
rect 531378 208350 531998 225922
rect 556590 226350 557066 226384
rect 556590 226294 556614 226350
rect 556670 226294 556738 226350
rect 556794 226294 556862 226350
rect 556918 226294 556986 226350
rect 557042 226294 557066 226350
rect 556590 226226 557066 226294
rect 556590 226170 556614 226226
rect 556670 226170 556738 226226
rect 556794 226170 556862 226226
rect 556918 226170 556986 226226
rect 557042 226170 557066 226226
rect 556590 226102 557066 226170
rect 556590 226046 556614 226102
rect 556670 226046 556738 226102
rect 556794 226046 556862 226102
rect 556918 226046 556986 226102
rect 557042 226046 557066 226102
rect 556590 225978 557066 226046
rect 556590 225922 556614 225978
rect 556670 225922 556738 225978
rect 556794 225922 556862 225978
rect 556918 225922 556986 225978
rect 557042 225922 557066 225978
rect 556590 225888 557066 225922
rect 557390 220350 557866 220384
rect 557390 220294 557414 220350
rect 557470 220294 557538 220350
rect 557594 220294 557662 220350
rect 557718 220294 557786 220350
rect 557842 220294 557866 220350
rect 557390 220226 557866 220294
rect 557390 220170 557414 220226
rect 557470 220170 557538 220226
rect 557594 220170 557662 220226
rect 557718 220170 557786 220226
rect 557842 220170 557866 220226
rect 557390 220102 557866 220170
rect 557390 220046 557414 220102
rect 557470 220046 557538 220102
rect 557594 220046 557662 220102
rect 557718 220046 557786 220102
rect 557842 220046 557866 220102
rect 557390 219978 557866 220046
rect 557390 219922 557414 219978
rect 557470 219922 557538 219978
rect 557594 219922 557662 219978
rect 557718 219922 557786 219978
rect 557842 219922 557866 219978
rect 557390 219888 557866 219922
rect 558378 220350 558998 237922
rect 558378 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 558998 220350
rect 558378 220226 558998 220294
rect 558378 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 558998 220226
rect 558378 220102 558998 220170
rect 558378 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 558998 220102
rect 558378 219978 558998 220046
rect 558378 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 558998 219978
rect 531378 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 531998 208350
rect 531378 208226 531998 208294
rect 531378 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 531998 208226
rect 531378 208102 531998 208170
rect 531378 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 531998 208102
rect 531378 207978 531998 208046
rect 531378 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 531998 207978
rect 531378 190350 531998 207922
rect 556590 208350 557066 208384
rect 556590 208294 556614 208350
rect 556670 208294 556738 208350
rect 556794 208294 556862 208350
rect 556918 208294 556986 208350
rect 557042 208294 557066 208350
rect 556590 208226 557066 208294
rect 556590 208170 556614 208226
rect 556670 208170 556738 208226
rect 556794 208170 556862 208226
rect 556918 208170 556986 208226
rect 557042 208170 557066 208226
rect 556590 208102 557066 208170
rect 556590 208046 556614 208102
rect 556670 208046 556738 208102
rect 556794 208046 556862 208102
rect 556918 208046 556986 208102
rect 557042 208046 557066 208102
rect 556590 207978 557066 208046
rect 556590 207922 556614 207978
rect 556670 207922 556738 207978
rect 556794 207922 556862 207978
rect 556918 207922 556986 207978
rect 557042 207922 557066 207978
rect 556590 207888 557066 207922
rect 557390 202350 557866 202384
rect 557390 202294 557414 202350
rect 557470 202294 557538 202350
rect 557594 202294 557662 202350
rect 557718 202294 557786 202350
rect 557842 202294 557866 202350
rect 557390 202226 557866 202294
rect 557390 202170 557414 202226
rect 557470 202170 557538 202226
rect 557594 202170 557662 202226
rect 557718 202170 557786 202226
rect 557842 202170 557866 202226
rect 557390 202102 557866 202170
rect 557390 202046 557414 202102
rect 557470 202046 557538 202102
rect 557594 202046 557662 202102
rect 557718 202046 557786 202102
rect 557842 202046 557866 202102
rect 557390 201978 557866 202046
rect 557390 201922 557414 201978
rect 557470 201922 557538 201978
rect 557594 201922 557662 201978
rect 557718 201922 557786 201978
rect 557842 201922 557866 201978
rect 557390 201888 557866 201922
rect 558378 202350 558998 219922
rect 558378 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 558998 202350
rect 558378 202226 558998 202294
rect 558378 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 558998 202226
rect 558378 202102 558998 202170
rect 558378 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 558998 202102
rect 558378 201978 558998 202046
rect 558378 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 558998 201978
rect 531378 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 531998 190350
rect 531378 190226 531998 190294
rect 531378 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 531998 190226
rect 531378 190102 531998 190170
rect 531378 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 531998 190102
rect 531378 189978 531998 190046
rect 531378 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 531998 189978
rect 531378 172350 531998 189922
rect 556590 190350 557066 190384
rect 556590 190294 556614 190350
rect 556670 190294 556738 190350
rect 556794 190294 556862 190350
rect 556918 190294 556986 190350
rect 557042 190294 557066 190350
rect 556590 190226 557066 190294
rect 556590 190170 556614 190226
rect 556670 190170 556738 190226
rect 556794 190170 556862 190226
rect 556918 190170 556986 190226
rect 557042 190170 557066 190226
rect 556590 190102 557066 190170
rect 556590 190046 556614 190102
rect 556670 190046 556738 190102
rect 556794 190046 556862 190102
rect 556918 190046 556986 190102
rect 557042 190046 557066 190102
rect 556590 189978 557066 190046
rect 556590 189922 556614 189978
rect 556670 189922 556738 189978
rect 556794 189922 556862 189978
rect 556918 189922 556986 189978
rect 557042 189922 557066 189978
rect 556590 189888 557066 189922
rect 557390 184350 557866 184384
rect 557390 184294 557414 184350
rect 557470 184294 557538 184350
rect 557594 184294 557662 184350
rect 557718 184294 557786 184350
rect 557842 184294 557866 184350
rect 557390 184226 557866 184294
rect 557390 184170 557414 184226
rect 557470 184170 557538 184226
rect 557594 184170 557662 184226
rect 557718 184170 557786 184226
rect 557842 184170 557866 184226
rect 557390 184102 557866 184170
rect 557390 184046 557414 184102
rect 557470 184046 557538 184102
rect 557594 184046 557662 184102
rect 557718 184046 557786 184102
rect 557842 184046 557866 184102
rect 557390 183978 557866 184046
rect 557390 183922 557414 183978
rect 557470 183922 557538 183978
rect 557594 183922 557662 183978
rect 557718 183922 557786 183978
rect 557842 183922 557866 183978
rect 557390 183888 557866 183922
rect 558378 184350 558998 201922
rect 558378 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 558998 184350
rect 558378 184226 558998 184294
rect 558378 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 558998 184226
rect 558378 184102 558998 184170
rect 558378 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 558998 184102
rect 558378 183978 558998 184046
rect 558378 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 558998 183978
rect 531378 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 531998 172350
rect 531378 172226 531998 172294
rect 531378 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 531998 172226
rect 531378 172102 531998 172170
rect 531378 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 531998 172102
rect 531378 171978 531998 172046
rect 531378 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 531998 171978
rect 531378 154350 531998 171922
rect 556590 172350 557066 172384
rect 556590 172294 556614 172350
rect 556670 172294 556738 172350
rect 556794 172294 556862 172350
rect 556918 172294 556986 172350
rect 557042 172294 557066 172350
rect 556590 172226 557066 172294
rect 556590 172170 556614 172226
rect 556670 172170 556738 172226
rect 556794 172170 556862 172226
rect 556918 172170 556986 172226
rect 557042 172170 557066 172226
rect 556590 172102 557066 172170
rect 556590 172046 556614 172102
rect 556670 172046 556738 172102
rect 556794 172046 556862 172102
rect 556918 172046 556986 172102
rect 557042 172046 557066 172102
rect 556590 171978 557066 172046
rect 556590 171922 556614 171978
rect 556670 171922 556738 171978
rect 556794 171922 556862 171978
rect 556918 171922 556986 171978
rect 557042 171922 557066 171978
rect 556590 171888 557066 171922
rect 557390 166350 557866 166384
rect 557390 166294 557414 166350
rect 557470 166294 557538 166350
rect 557594 166294 557662 166350
rect 557718 166294 557786 166350
rect 557842 166294 557866 166350
rect 557390 166226 557866 166294
rect 557390 166170 557414 166226
rect 557470 166170 557538 166226
rect 557594 166170 557662 166226
rect 557718 166170 557786 166226
rect 557842 166170 557866 166226
rect 557390 166102 557866 166170
rect 557390 166046 557414 166102
rect 557470 166046 557538 166102
rect 557594 166046 557662 166102
rect 557718 166046 557786 166102
rect 557842 166046 557866 166102
rect 557390 165978 557866 166046
rect 557390 165922 557414 165978
rect 557470 165922 557538 165978
rect 557594 165922 557662 165978
rect 557718 165922 557786 165978
rect 557842 165922 557866 165978
rect 557390 165888 557866 165922
rect 558378 166350 558998 183922
rect 558378 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 558998 166350
rect 558378 166226 558998 166294
rect 558378 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 558998 166226
rect 558378 166102 558998 166170
rect 558378 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 558998 166102
rect 558378 165978 558998 166046
rect 558378 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 558998 165978
rect 531378 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 531998 154350
rect 531378 154226 531998 154294
rect 531378 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 531998 154226
rect 531378 154102 531998 154170
rect 531378 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 531998 154102
rect 531378 153978 531998 154046
rect 531378 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 531998 153978
rect 531378 136350 531998 153922
rect 558378 148350 558998 165922
rect 558378 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 558998 148350
rect 558378 148226 558998 148294
rect 558378 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 558998 148226
rect 558378 148102 558998 148170
rect 558378 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 558998 148102
rect 558378 147978 558998 148046
rect 558378 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 558998 147978
rect 544684 142498 544740 142508
rect 534604 141958 534660 141968
rect 534604 141204 534660 141902
rect 534604 141138 534660 141148
rect 544684 141204 544740 142442
rect 544684 141138 544740 141148
rect 531378 136294 531474 136350
rect 531530 136294 531598 136350
rect 531654 136294 531722 136350
rect 531778 136294 531846 136350
rect 531902 136294 531998 136350
rect 531378 136226 531998 136294
rect 531378 136170 531474 136226
rect 531530 136170 531598 136226
rect 531654 136170 531722 136226
rect 531778 136170 531846 136226
rect 531902 136170 531998 136226
rect 531378 136102 531998 136170
rect 531378 136046 531474 136102
rect 531530 136046 531598 136102
rect 531654 136046 531722 136102
rect 531778 136046 531846 136102
rect 531902 136046 531998 136102
rect 531378 135978 531998 136046
rect 531378 135922 531474 135978
rect 531530 135922 531598 135978
rect 531654 135922 531722 135978
rect 531778 135922 531846 135978
rect 531902 135922 531998 135978
rect 531378 118350 531998 135922
rect 545788 130350 546264 130384
rect 545788 130294 545812 130350
rect 545868 130294 545936 130350
rect 545992 130294 546060 130350
rect 546116 130294 546184 130350
rect 546240 130294 546264 130350
rect 545788 130226 546264 130294
rect 545788 130170 545812 130226
rect 545868 130170 545936 130226
rect 545992 130170 546060 130226
rect 546116 130170 546184 130226
rect 546240 130170 546264 130226
rect 545788 130102 546264 130170
rect 545788 130046 545812 130102
rect 545868 130046 545936 130102
rect 545992 130046 546060 130102
rect 546116 130046 546184 130102
rect 546240 130046 546264 130102
rect 545788 129978 546264 130046
rect 545788 129922 545812 129978
rect 545868 129922 545936 129978
rect 545992 129922 546060 129978
rect 546116 129922 546184 129978
rect 546240 129922 546264 129978
rect 545788 129888 546264 129922
rect 558378 130350 558998 147922
rect 558378 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 558998 130350
rect 558378 130226 558998 130294
rect 558378 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 558998 130226
rect 558378 130102 558998 130170
rect 558378 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 558998 130102
rect 558378 129978 558998 130046
rect 558378 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 558998 129978
rect 531378 118294 531474 118350
rect 531530 118294 531598 118350
rect 531654 118294 531722 118350
rect 531778 118294 531846 118350
rect 531902 118294 531998 118350
rect 531378 118226 531998 118294
rect 531378 118170 531474 118226
rect 531530 118170 531598 118226
rect 531654 118170 531722 118226
rect 531778 118170 531846 118226
rect 531902 118170 531998 118226
rect 531378 118102 531998 118170
rect 531378 118046 531474 118102
rect 531530 118046 531598 118102
rect 531654 118046 531722 118102
rect 531778 118046 531846 118102
rect 531902 118046 531998 118102
rect 531378 117978 531998 118046
rect 531378 117922 531474 117978
rect 531530 117922 531598 117978
rect 531654 117922 531722 117978
rect 531778 117922 531846 117978
rect 531902 117922 531998 117978
rect 531378 100350 531998 117922
rect 546588 118350 547064 118384
rect 546588 118294 546612 118350
rect 546668 118294 546736 118350
rect 546792 118294 546860 118350
rect 546916 118294 546984 118350
rect 547040 118294 547064 118350
rect 546588 118226 547064 118294
rect 546588 118170 546612 118226
rect 546668 118170 546736 118226
rect 546792 118170 546860 118226
rect 546916 118170 546984 118226
rect 547040 118170 547064 118226
rect 546588 118102 547064 118170
rect 546588 118046 546612 118102
rect 546668 118046 546736 118102
rect 546792 118046 546860 118102
rect 546916 118046 546984 118102
rect 547040 118046 547064 118102
rect 546588 117978 547064 118046
rect 546588 117922 546612 117978
rect 546668 117922 546736 117978
rect 546792 117922 546860 117978
rect 546916 117922 546984 117978
rect 547040 117922 547064 117978
rect 546588 117888 547064 117922
rect 545788 112350 546264 112384
rect 545788 112294 545812 112350
rect 545868 112294 545936 112350
rect 545992 112294 546060 112350
rect 546116 112294 546184 112350
rect 546240 112294 546264 112350
rect 545788 112226 546264 112294
rect 545788 112170 545812 112226
rect 545868 112170 545936 112226
rect 545992 112170 546060 112226
rect 546116 112170 546184 112226
rect 546240 112170 546264 112226
rect 545788 112102 546264 112170
rect 545788 112046 545812 112102
rect 545868 112046 545936 112102
rect 545992 112046 546060 112102
rect 546116 112046 546184 112102
rect 546240 112046 546264 112102
rect 545788 111978 546264 112046
rect 545788 111922 545812 111978
rect 545868 111922 545936 111978
rect 545992 111922 546060 111978
rect 546116 111922 546184 111978
rect 546240 111922 546264 111978
rect 545788 111888 546264 111922
rect 558378 112350 558998 129922
rect 558378 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 558998 112350
rect 558378 112226 558998 112294
rect 558378 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 558998 112226
rect 558378 112102 558998 112170
rect 558378 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 558998 112102
rect 558378 111978 558998 112046
rect 558378 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 558998 111978
rect 531378 100294 531474 100350
rect 531530 100294 531598 100350
rect 531654 100294 531722 100350
rect 531778 100294 531846 100350
rect 531902 100294 531998 100350
rect 531378 100226 531998 100294
rect 531378 100170 531474 100226
rect 531530 100170 531598 100226
rect 531654 100170 531722 100226
rect 531778 100170 531846 100226
rect 531902 100170 531998 100226
rect 531378 100102 531998 100170
rect 531378 100046 531474 100102
rect 531530 100046 531598 100102
rect 531654 100046 531722 100102
rect 531778 100046 531846 100102
rect 531902 100046 531998 100102
rect 531378 99978 531998 100046
rect 531378 99922 531474 99978
rect 531530 99922 531598 99978
rect 531654 99922 531722 99978
rect 531778 99922 531846 99978
rect 531902 99922 531998 99978
rect 531378 82350 531998 99922
rect 546588 100350 547064 100384
rect 546588 100294 546612 100350
rect 546668 100294 546736 100350
rect 546792 100294 546860 100350
rect 546916 100294 546984 100350
rect 547040 100294 547064 100350
rect 546588 100226 547064 100294
rect 546588 100170 546612 100226
rect 546668 100170 546736 100226
rect 546792 100170 546860 100226
rect 546916 100170 546984 100226
rect 547040 100170 547064 100226
rect 546588 100102 547064 100170
rect 546588 100046 546612 100102
rect 546668 100046 546736 100102
rect 546792 100046 546860 100102
rect 546916 100046 546984 100102
rect 547040 100046 547064 100102
rect 546588 99978 547064 100046
rect 546588 99922 546612 99978
rect 546668 99922 546736 99978
rect 546792 99922 546860 99978
rect 546916 99922 546984 99978
rect 547040 99922 547064 99978
rect 546588 99888 547064 99922
rect 545788 94350 546264 94384
rect 545788 94294 545812 94350
rect 545868 94294 545936 94350
rect 545992 94294 546060 94350
rect 546116 94294 546184 94350
rect 546240 94294 546264 94350
rect 545788 94226 546264 94294
rect 545788 94170 545812 94226
rect 545868 94170 545936 94226
rect 545992 94170 546060 94226
rect 546116 94170 546184 94226
rect 546240 94170 546264 94226
rect 545788 94102 546264 94170
rect 545788 94046 545812 94102
rect 545868 94046 545936 94102
rect 545992 94046 546060 94102
rect 546116 94046 546184 94102
rect 546240 94046 546264 94102
rect 545788 93978 546264 94046
rect 545788 93922 545812 93978
rect 545868 93922 545936 93978
rect 545992 93922 546060 93978
rect 546116 93922 546184 93978
rect 546240 93922 546264 93978
rect 545788 93888 546264 93922
rect 558378 94350 558998 111922
rect 558378 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 558998 94350
rect 558378 94226 558998 94294
rect 558378 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 558998 94226
rect 558378 94102 558998 94170
rect 558378 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 558998 94102
rect 558378 93978 558998 94046
rect 558378 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 558998 93978
rect 531378 82294 531474 82350
rect 531530 82294 531598 82350
rect 531654 82294 531722 82350
rect 531778 82294 531846 82350
rect 531902 82294 531998 82350
rect 531378 82226 531998 82294
rect 531378 82170 531474 82226
rect 531530 82170 531598 82226
rect 531654 82170 531722 82226
rect 531778 82170 531846 82226
rect 531902 82170 531998 82226
rect 531378 82102 531998 82170
rect 531378 82046 531474 82102
rect 531530 82046 531598 82102
rect 531654 82046 531722 82102
rect 531778 82046 531846 82102
rect 531902 82046 531998 82102
rect 531378 81978 531998 82046
rect 531378 81922 531474 81978
rect 531530 81922 531598 81978
rect 531654 81922 531722 81978
rect 531778 81922 531846 81978
rect 531902 81922 531998 81978
rect 531378 64350 531998 81922
rect 546588 82350 547064 82384
rect 546588 82294 546612 82350
rect 546668 82294 546736 82350
rect 546792 82294 546860 82350
rect 546916 82294 546984 82350
rect 547040 82294 547064 82350
rect 546588 82226 547064 82294
rect 546588 82170 546612 82226
rect 546668 82170 546736 82226
rect 546792 82170 546860 82226
rect 546916 82170 546984 82226
rect 547040 82170 547064 82226
rect 546588 82102 547064 82170
rect 546588 82046 546612 82102
rect 546668 82046 546736 82102
rect 546792 82046 546860 82102
rect 546916 82046 546984 82102
rect 547040 82046 547064 82102
rect 546588 81978 547064 82046
rect 546588 81922 546612 81978
rect 546668 81922 546736 81978
rect 546792 81922 546860 81978
rect 546916 81922 546984 81978
rect 547040 81922 547064 81978
rect 546588 81888 547064 81922
rect 545788 76350 546264 76384
rect 545788 76294 545812 76350
rect 545868 76294 545936 76350
rect 545992 76294 546060 76350
rect 546116 76294 546184 76350
rect 546240 76294 546264 76350
rect 545788 76226 546264 76294
rect 545788 76170 545812 76226
rect 545868 76170 545936 76226
rect 545992 76170 546060 76226
rect 546116 76170 546184 76226
rect 546240 76170 546264 76226
rect 545788 76102 546264 76170
rect 545788 76046 545812 76102
rect 545868 76046 545936 76102
rect 545992 76046 546060 76102
rect 546116 76046 546184 76102
rect 546240 76046 546264 76102
rect 545788 75978 546264 76046
rect 545788 75922 545812 75978
rect 545868 75922 545936 75978
rect 545992 75922 546060 75978
rect 546116 75922 546184 75978
rect 546240 75922 546264 75978
rect 545788 75888 546264 75922
rect 558378 76350 558998 93922
rect 558378 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 558998 76350
rect 558378 76226 558998 76294
rect 558378 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 558998 76226
rect 558378 76102 558998 76170
rect 558378 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 558998 76102
rect 558378 75978 558998 76046
rect 558378 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 558998 75978
rect 531378 64294 531474 64350
rect 531530 64294 531598 64350
rect 531654 64294 531722 64350
rect 531778 64294 531846 64350
rect 531902 64294 531998 64350
rect 531378 64226 531998 64294
rect 531378 64170 531474 64226
rect 531530 64170 531598 64226
rect 531654 64170 531722 64226
rect 531778 64170 531846 64226
rect 531902 64170 531998 64226
rect 531378 64102 531998 64170
rect 531378 64046 531474 64102
rect 531530 64046 531598 64102
rect 531654 64046 531722 64102
rect 531778 64046 531846 64102
rect 531902 64046 531998 64102
rect 531378 63978 531998 64046
rect 531378 63922 531474 63978
rect 531530 63922 531598 63978
rect 531654 63922 531722 63978
rect 531778 63922 531846 63978
rect 531902 63922 531998 63978
rect 531378 46350 531998 63922
rect 546588 64350 547064 64384
rect 546588 64294 546612 64350
rect 546668 64294 546736 64350
rect 546792 64294 546860 64350
rect 546916 64294 546984 64350
rect 547040 64294 547064 64350
rect 546588 64226 547064 64294
rect 546588 64170 546612 64226
rect 546668 64170 546736 64226
rect 546792 64170 546860 64226
rect 546916 64170 546984 64226
rect 547040 64170 547064 64226
rect 546588 64102 547064 64170
rect 546588 64046 546612 64102
rect 546668 64046 546736 64102
rect 546792 64046 546860 64102
rect 546916 64046 546984 64102
rect 547040 64046 547064 64102
rect 546588 63978 547064 64046
rect 546588 63922 546612 63978
rect 546668 63922 546736 63978
rect 546792 63922 546860 63978
rect 546916 63922 546984 63978
rect 547040 63922 547064 63978
rect 546588 63888 547064 63922
rect 545788 58350 546264 58384
rect 545788 58294 545812 58350
rect 545868 58294 545936 58350
rect 545992 58294 546060 58350
rect 546116 58294 546184 58350
rect 546240 58294 546264 58350
rect 545788 58226 546264 58294
rect 545788 58170 545812 58226
rect 545868 58170 545936 58226
rect 545992 58170 546060 58226
rect 546116 58170 546184 58226
rect 546240 58170 546264 58226
rect 545788 58102 546264 58170
rect 545788 58046 545812 58102
rect 545868 58046 545936 58102
rect 545992 58046 546060 58102
rect 546116 58046 546184 58102
rect 546240 58046 546264 58102
rect 545788 57978 546264 58046
rect 545788 57922 545812 57978
rect 545868 57922 545936 57978
rect 545992 57922 546060 57978
rect 546116 57922 546184 57978
rect 546240 57922 546264 57978
rect 545788 57888 546264 57922
rect 558378 58350 558998 75922
rect 558378 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 558998 58350
rect 558378 58226 558998 58294
rect 558378 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 558998 58226
rect 558378 58102 558998 58170
rect 558378 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 558998 58102
rect 558378 57978 558998 58046
rect 558378 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 558998 57978
rect 531378 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 531998 46350
rect 531378 46226 531998 46294
rect 531378 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 531998 46226
rect 531378 46102 531998 46170
rect 531378 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 531998 46102
rect 531378 45978 531998 46046
rect 531378 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 531998 45978
rect 531378 28350 531998 45922
rect 546588 46350 547064 46384
rect 546588 46294 546612 46350
rect 546668 46294 546736 46350
rect 546792 46294 546860 46350
rect 546916 46294 546984 46350
rect 547040 46294 547064 46350
rect 546588 46226 547064 46294
rect 546588 46170 546612 46226
rect 546668 46170 546736 46226
rect 546792 46170 546860 46226
rect 546916 46170 546984 46226
rect 547040 46170 547064 46226
rect 546588 46102 547064 46170
rect 546588 46046 546612 46102
rect 546668 46046 546736 46102
rect 546792 46046 546860 46102
rect 546916 46046 546984 46102
rect 547040 46046 547064 46102
rect 546588 45978 547064 46046
rect 546588 45922 546612 45978
rect 546668 45922 546736 45978
rect 546792 45922 546860 45978
rect 546916 45922 546984 45978
rect 547040 45922 547064 45978
rect 546588 45888 547064 45922
rect 531378 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 531998 28350
rect 531378 28226 531998 28294
rect 531378 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 531998 28226
rect 531378 28102 531998 28170
rect 531378 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 531998 28102
rect 531378 27978 531998 28046
rect 531378 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 531998 27978
rect 531378 10350 531998 27922
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 531378 -1120 531998 9922
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 40350 558998 57922
rect 558378 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 558998 40350
rect 558378 40226 558998 40294
rect 558378 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 558998 40226
rect 558378 40102 558998 40170
rect 558378 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 558998 40102
rect 558378 39978 558998 40046
rect 558378 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 558998 39978
rect 558378 22350 558998 39922
rect 558378 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 558998 22350
rect 558378 22226 558998 22294
rect 558378 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 558998 22226
rect 558378 22102 558998 22170
rect 558378 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 558998 22102
rect 558378 21978 558998 22046
rect 558378 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 558998 21978
rect 558378 4350 558998 21922
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 558378 -160 558998 3922
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 584668 591332 584724 591342
rect 584668 589798 584724 591276
rect 584668 589732 584724 589742
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 562098 550350 562718 567922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 562098 532350 562718 549922
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 562098 478350 562718 495922
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 562098 460350 562718 477922
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 562098 388350 562718 405922
rect 562098 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 562718 388350
rect 562098 388226 562718 388294
rect 562098 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 562718 388226
rect 562098 388102 562718 388170
rect 562098 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 562718 388102
rect 562098 387978 562718 388046
rect 562098 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 562718 387978
rect 562098 370350 562718 387922
rect 562098 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 562718 370350
rect 562098 370226 562718 370294
rect 562098 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 562718 370226
rect 562098 370102 562718 370170
rect 562098 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 562718 370102
rect 562098 369978 562718 370046
rect 562098 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 562718 369978
rect 562098 352350 562718 369922
rect 562098 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 562718 352350
rect 562098 352226 562718 352294
rect 562098 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 562718 352226
rect 562098 352102 562718 352170
rect 562098 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 562718 352102
rect 562098 351978 562718 352046
rect 562098 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 562718 351978
rect 562098 334350 562718 351922
rect 562098 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 562718 334350
rect 562098 334226 562718 334294
rect 562098 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 562718 334226
rect 562098 334102 562718 334170
rect 562098 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 562718 334102
rect 562098 333978 562718 334046
rect 562098 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 562718 333978
rect 562098 316350 562718 333922
rect 562098 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 562718 316350
rect 562098 316226 562718 316294
rect 562098 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 562718 316226
rect 562098 316102 562718 316170
rect 562098 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 562718 316102
rect 562098 315978 562718 316046
rect 562098 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 562718 315978
rect 562098 298350 562718 315922
rect 562098 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 562718 298350
rect 562098 298226 562718 298294
rect 562098 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 562718 298226
rect 562098 298102 562718 298170
rect 562098 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 562718 298102
rect 562098 297978 562718 298046
rect 562098 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 562718 297978
rect 562098 280350 562718 297922
rect 562098 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 562718 280350
rect 562098 280226 562718 280294
rect 562098 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 562718 280226
rect 562098 280102 562718 280170
rect 562098 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 562718 280102
rect 562098 279978 562718 280046
rect 562098 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 562718 279978
rect 562098 262350 562718 279922
rect 589098 580350 589718 596784
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 589098 562350 589718 579922
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 590604 551098 590660 551108
rect 590156 548996 590212 549006
rect 590156 547858 590212 548940
rect 590156 547792 590212 547802
rect 590492 548038 590548 548048
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 590492 522788 590548 547982
rect 590604 535892 590660 551042
rect 590604 535826 590660 535836
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 590492 522722 590548 522732
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 590716 509348 590772 509358
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 589098 400350 589718 417922
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 589098 382350 589718 399922
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 589098 364350 589718 381922
rect 590492 496132 590548 496142
rect 590156 377188 590212 377198
rect 590156 376498 590212 377132
rect 590156 376432 590212 376442
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 589098 292350 589718 309922
rect 590492 295498 590548 496076
rect 590492 295432 590548 295442
rect 590604 456484 590660 456494
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 589098 274350 589718 291922
rect 590156 285238 590212 285248
rect 590156 284900 590212 285182
rect 590156 284834 590212 284844
rect 590604 281998 590660 456428
rect 590716 451018 590772 509292
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 590716 450952 590772 450962
rect 590828 469700 590884 469710
rect 590828 450660 590884 469644
rect 590828 450594 590884 450604
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 590828 430164 590884 430174
rect 590716 416836 590772 416846
rect 590716 285598 590772 416780
rect 590828 301618 590884 430108
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 591052 403620 591108 403630
rect 590828 301552 590884 301562
rect 590940 390404 590996 390414
rect 590940 300718 590996 390348
rect 591052 387658 591108 403564
rect 591052 387592 591108 387602
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 590940 300652 590996 300662
rect 591052 350756 591108 350766
rect 590716 285532 590772 285542
rect 590828 297892 590884 297902
rect 590828 282178 590884 297836
rect 591052 297298 591108 350700
rect 591052 297232 591108 297242
rect 591164 337540 591220 337550
rect 591164 288838 591220 337484
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 591276 311108 591332 311118
rect 591276 295678 591332 311052
rect 591276 295612 591332 295622
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 591164 288772 591220 288782
rect 590828 282112 590884 282122
rect 590604 281932 590660 281942
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 562098 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 562718 262350
rect 562098 262226 562718 262294
rect 562098 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 562718 262226
rect 562098 262102 562718 262170
rect 562098 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 562718 262102
rect 562098 261978 562718 262046
rect 562098 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 562718 261978
rect 562098 244350 562718 261922
rect 562098 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 562718 244350
rect 562098 244226 562718 244294
rect 562098 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 562718 244226
rect 562098 244102 562718 244170
rect 562098 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 562718 244102
rect 562098 243978 562718 244046
rect 562098 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 562718 243978
rect 562098 226350 562718 243922
rect 562098 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 562718 226350
rect 562098 226226 562718 226294
rect 562098 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 562718 226226
rect 562098 226102 562718 226170
rect 562098 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 562718 226102
rect 562098 225978 562718 226046
rect 562098 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 562718 225978
rect 562098 208350 562718 225922
rect 562098 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 562718 208350
rect 562098 208226 562718 208294
rect 562098 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 562718 208226
rect 562098 208102 562718 208170
rect 562098 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 562718 208102
rect 562098 207978 562718 208046
rect 562098 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 562718 207978
rect 562098 190350 562718 207922
rect 562098 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 562718 190350
rect 562098 190226 562718 190294
rect 562098 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 562718 190226
rect 562098 190102 562718 190170
rect 562098 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 562718 190102
rect 562098 189978 562718 190046
rect 562098 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 562718 189978
rect 562098 172350 562718 189922
rect 562098 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 562718 172350
rect 562098 172226 562718 172294
rect 562098 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 562718 172226
rect 562098 172102 562718 172170
rect 562098 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 562718 172102
rect 562098 171978 562718 172046
rect 562098 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 562718 171978
rect 562098 154350 562718 171922
rect 562098 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 562718 154350
rect 562098 154226 562718 154294
rect 562098 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 562718 154226
rect 562098 154102 562718 154170
rect 562098 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 562718 154102
rect 562098 153978 562718 154046
rect 562098 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 562718 153978
rect 562098 136350 562718 153922
rect 562098 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 562718 136350
rect 562098 136226 562718 136294
rect 562098 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 562718 136226
rect 562098 136102 562718 136170
rect 562098 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 562718 136102
rect 562098 135978 562718 136046
rect 562098 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 562718 135978
rect 562098 118350 562718 135922
rect 562098 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 562718 118350
rect 562098 118226 562718 118294
rect 562098 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 562718 118226
rect 562098 118102 562718 118170
rect 562098 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 562718 118102
rect 562098 117978 562718 118046
rect 562098 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 562718 117978
rect 562098 100350 562718 117922
rect 562098 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 562718 100350
rect 562098 100226 562718 100294
rect 562098 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 562718 100226
rect 562098 100102 562718 100170
rect 562098 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 562718 100102
rect 562098 99978 562718 100046
rect 562098 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 562718 99978
rect 562098 82350 562718 99922
rect 562098 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 562718 82350
rect 562098 82226 562718 82294
rect 562098 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 562718 82226
rect 562098 82102 562718 82170
rect 562098 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 562718 82102
rect 562098 81978 562718 82046
rect 562098 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 562718 81978
rect 562098 64350 562718 81922
rect 562098 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 562718 64350
rect 562098 64226 562718 64294
rect 562098 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 562718 64226
rect 562098 64102 562718 64170
rect 562098 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 562718 64102
rect 562098 63978 562718 64046
rect 562098 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 562718 63978
rect 562098 46350 562718 63922
rect 566972 271348 567028 271358
rect 566972 60004 567028 271292
rect 572012 267988 572068 267998
rect 572012 258244 572068 267932
rect 572012 258178 572068 258188
rect 566972 59938 567028 59948
rect 589098 256350 589718 273922
rect 590828 278068 590884 278078
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 589098 238350 589718 255922
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 590492 273028 590548 273038
rect 590156 206398 590212 206408
rect 590156 205604 590212 206342
rect 590156 205538 590212 205548
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 589098 148350 589718 165922
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 589098 130350 589718 147922
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 590156 127558 590212 127568
rect 590156 126308 590212 127502
rect 590156 126242 590212 126252
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 589098 94350 589718 111922
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 589098 76350 589718 93922
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 562098 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 562718 46350
rect 562098 46226 562718 46294
rect 562098 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 562718 46226
rect 562098 46102 562718 46170
rect 562098 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 562718 46102
rect 562098 45978 562718 46046
rect 562098 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 562718 45978
rect 562098 28350 562718 45922
rect 562098 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 562718 28350
rect 562098 28226 562718 28294
rect 562098 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 562718 28226
rect 562098 28102 562718 28170
rect 562098 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 562718 28102
rect 562098 27978 562718 28046
rect 562098 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 562718 27978
rect 562098 10350 562718 27922
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 562098 -1120 562718 9922
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 58350 589718 75922
rect 590492 73444 590548 272972
rect 590716 261268 590772 261278
rect 590604 259588 590660 259598
rect 590604 192388 590660 259532
rect 590716 218820 590772 261212
rect 590828 232036 590884 278012
rect 590828 231970 590884 231980
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 590716 218754 590772 218764
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 590604 192322 590660 192332
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 590828 160580 590884 160590
rect 590604 145348 590660 145358
rect 590604 113092 590660 145292
rect 590604 113026 590660 113036
rect 590828 99876 590884 160524
rect 590828 99810 590884 99820
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 590492 73378 590548 73388
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 589098 40350 589718 57922
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 589098 22350 589718 39922
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 589098 4350 589718 21922
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect 4172 557882 4228 557938
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect 4172 551222 4228 551278
rect 4284 548162 4340 548218
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 4956 430802 5012 430858
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect 4172 430082 4228 430138
rect 4284 426842 4340 426898
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect 4172 347642 4228 347698
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect 4172 300482 4228 300538
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect 4284 293822 4340 293878
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 4396 288602 4452 288658
rect 4956 283742 5012 283798
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 4172 248500 4228 248518
rect 4172 248462 4228 248500
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 4172 235142 4228 235198
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect 4172 206522 4228 206578
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 9234 370294 9290 370350
rect 9358 370294 9414 370350
rect 9482 370294 9538 370350
rect 9606 370294 9662 370350
rect 9234 370170 9290 370226
rect 9358 370170 9414 370226
rect 9482 370170 9538 370226
rect 9606 370170 9662 370226
rect 9234 370046 9290 370102
rect 9358 370046 9414 370102
rect 9482 370046 9538 370102
rect 9606 370046 9662 370102
rect 9234 369922 9290 369978
rect 9358 369922 9414 369978
rect 9482 369922 9538 369978
rect 9606 369922 9662 369978
rect 9234 352294 9290 352350
rect 9358 352294 9414 352350
rect 9482 352294 9538 352350
rect 9606 352294 9662 352350
rect 9234 352170 9290 352226
rect 9358 352170 9414 352226
rect 9482 352170 9538 352226
rect 9606 352170 9662 352226
rect 9234 352046 9290 352102
rect 9358 352046 9414 352102
rect 9482 352046 9538 352102
rect 9606 352046 9662 352102
rect 9234 351922 9290 351978
rect 9358 351922 9414 351978
rect 9482 351922 9538 351978
rect 9606 351922 9662 351978
rect 9234 334294 9290 334350
rect 9358 334294 9414 334350
rect 9482 334294 9538 334350
rect 9606 334294 9662 334350
rect 9234 334170 9290 334226
rect 9358 334170 9414 334226
rect 9482 334170 9538 334226
rect 9606 334170 9662 334226
rect 9234 334046 9290 334102
rect 9358 334046 9414 334102
rect 9482 334046 9538 334102
rect 9606 334046 9662 334102
rect 9234 333922 9290 333978
rect 9358 333922 9414 333978
rect 9482 333922 9538 333978
rect 9606 333922 9662 333978
rect 9234 316294 9290 316350
rect 9358 316294 9414 316350
rect 9482 316294 9538 316350
rect 9606 316294 9662 316350
rect 9234 316170 9290 316226
rect 9358 316170 9414 316226
rect 9482 316170 9538 316226
rect 9606 316170 9662 316226
rect 9234 316046 9290 316102
rect 9358 316046 9414 316102
rect 9482 316046 9538 316102
rect 9606 316046 9662 316102
rect 9234 315922 9290 315978
rect 9358 315922 9414 315978
rect 9482 315922 9538 315978
rect 9606 315922 9662 315978
rect 9234 298294 9290 298350
rect 9358 298294 9414 298350
rect 9482 298294 9538 298350
rect 9606 298294 9662 298350
rect 9234 298170 9290 298226
rect 9358 298170 9414 298226
rect 9482 298170 9538 298226
rect 9606 298170 9662 298226
rect 9234 298046 9290 298102
rect 9358 298046 9414 298102
rect 9482 298046 9538 298102
rect 9606 298046 9662 298102
rect 9234 297922 9290 297978
rect 9358 297922 9414 297978
rect 9482 297922 9538 297978
rect 9606 297922 9662 297978
rect 9234 280294 9290 280350
rect 9358 280294 9414 280350
rect 9482 280294 9538 280350
rect 9606 280294 9662 280350
rect 9234 280170 9290 280226
rect 9358 280170 9414 280226
rect 9482 280170 9538 280226
rect 9606 280170 9662 280226
rect 9234 280046 9290 280102
rect 9358 280046 9414 280102
rect 9482 280046 9538 280102
rect 9606 280046 9662 280102
rect 9234 279922 9290 279978
rect 9358 279922 9414 279978
rect 9482 279922 9538 279978
rect 9606 279922 9662 279978
rect 9234 262294 9290 262350
rect 9358 262294 9414 262350
rect 9482 262294 9538 262350
rect 9606 262294 9662 262350
rect 9234 262170 9290 262226
rect 9358 262170 9414 262226
rect 9482 262170 9538 262226
rect 9606 262170 9662 262226
rect 9234 262046 9290 262102
rect 9358 262046 9414 262102
rect 9482 262046 9538 262102
rect 9606 262046 9662 262102
rect 9234 261922 9290 261978
rect 9358 261922 9414 261978
rect 9482 261922 9538 261978
rect 9606 261922 9662 261978
rect 9234 244294 9290 244350
rect 9358 244294 9414 244350
rect 9482 244294 9538 244350
rect 9606 244294 9662 244350
rect 9234 244170 9290 244226
rect 9358 244170 9414 244226
rect 9482 244170 9538 244226
rect 9606 244170 9662 244226
rect 9234 244046 9290 244102
rect 9358 244046 9414 244102
rect 9482 244046 9538 244102
rect 9606 244046 9662 244102
rect 9234 243922 9290 243978
rect 9358 243922 9414 243978
rect 9482 243922 9538 243978
rect 9606 243922 9662 243978
rect 9234 226294 9290 226350
rect 9358 226294 9414 226350
rect 9482 226294 9538 226350
rect 9606 226294 9662 226350
rect 9234 226170 9290 226226
rect 9358 226170 9414 226226
rect 9482 226170 9538 226226
rect 9606 226170 9662 226226
rect 9234 226046 9290 226102
rect 9358 226046 9414 226102
rect 9482 226046 9538 226102
rect 9606 226046 9662 226102
rect 9234 225922 9290 225978
rect 9358 225922 9414 225978
rect 9482 225922 9538 225978
rect 9606 225922 9662 225978
rect 9234 208294 9290 208350
rect 9358 208294 9414 208350
rect 9482 208294 9538 208350
rect 9606 208294 9662 208350
rect 9234 208170 9290 208226
rect 9358 208170 9414 208226
rect 9482 208170 9538 208226
rect 9606 208170 9662 208226
rect 9234 208046 9290 208102
rect 9358 208046 9414 208102
rect 9482 208046 9538 208102
rect 9606 208046 9662 208102
rect 9234 207922 9290 207978
rect 9358 207922 9414 207978
rect 9482 207922 9538 207978
rect 9606 207922 9662 207978
rect 9234 190294 9290 190350
rect 9358 190294 9414 190350
rect 9482 190294 9538 190350
rect 9606 190294 9662 190350
rect 9234 190170 9290 190226
rect 9358 190170 9414 190226
rect 9482 190170 9538 190226
rect 9606 190170 9662 190226
rect 9234 190046 9290 190102
rect 9358 190046 9414 190102
rect 9482 190046 9538 190102
rect 9606 190046 9662 190102
rect 9234 189922 9290 189978
rect 9358 189922 9414 189978
rect 9482 189922 9538 189978
rect 9606 189922 9662 189978
rect 9234 172294 9290 172350
rect 9358 172294 9414 172350
rect 9482 172294 9538 172350
rect 9606 172294 9662 172350
rect 9234 172170 9290 172226
rect 9358 172170 9414 172226
rect 9482 172170 9538 172226
rect 9606 172170 9662 172226
rect 9234 172046 9290 172102
rect 9358 172046 9414 172102
rect 9482 172046 9538 172102
rect 9606 172046 9662 172102
rect 9234 171922 9290 171978
rect 9358 171922 9414 171978
rect 9482 171922 9538 171978
rect 9606 171922 9662 171978
rect 9234 154294 9290 154350
rect 9358 154294 9414 154350
rect 9482 154294 9538 154350
rect 9606 154294 9662 154350
rect 9234 154170 9290 154226
rect 9358 154170 9414 154226
rect 9482 154170 9538 154226
rect 9606 154170 9662 154226
rect 9234 154046 9290 154102
rect 9358 154046 9414 154102
rect 9482 154046 9538 154102
rect 9606 154046 9662 154102
rect 9234 153922 9290 153978
rect 9358 153922 9414 153978
rect 9482 153922 9538 153978
rect 9606 153922 9662 153978
rect 9234 136294 9290 136350
rect 9358 136294 9414 136350
rect 9482 136294 9538 136350
rect 9606 136294 9662 136350
rect 9234 136170 9290 136226
rect 9358 136170 9414 136226
rect 9482 136170 9538 136226
rect 9606 136170 9662 136226
rect 9234 136046 9290 136102
rect 9358 136046 9414 136102
rect 9482 136046 9538 136102
rect 9606 136046 9662 136102
rect 9234 135922 9290 135978
rect 9358 135922 9414 135978
rect 9482 135922 9538 135978
rect 9606 135922 9662 135978
rect 9234 118294 9290 118350
rect 9358 118294 9414 118350
rect 9482 118294 9538 118350
rect 9606 118294 9662 118350
rect 9234 118170 9290 118226
rect 9358 118170 9414 118226
rect 9482 118170 9538 118226
rect 9606 118170 9662 118226
rect 9234 118046 9290 118102
rect 9358 118046 9414 118102
rect 9482 118046 9538 118102
rect 9606 118046 9662 118102
rect 9234 117922 9290 117978
rect 9358 117922 9414 117978
rect 9482 117922 9538 117978
rect 9606 117922 9662 117978
rect 9234 100294 9290 100350
rect 9358 100294 9414 100350
rect 9482 100294 9538 100350
rect 9606 100294 9662 100350
rect 9234 100170 9290 100226
rect 9358 100170 9414 100226
rect 9482 100170 9538 100226
rect 9606 100170 9662 100226
rect 9234 100046 9290 100102
rect 9358 100046 9414 100102
rect 9482 100046 9538 100102
rect 9606 100046 9662 100102
rect 9234 99922 9290 99978
rect 9358 99922 9414 99978
rect 9482 99922 9538 99978
rect 9606 99922 9662 99978
rect 9234 82294 9290 82350
rect 9358 82294 9414 82350
rect 9482 82294 9538 82350
rect 9606 82294 9662 82350
rect 9234 82170 9290 82226
rect 9358 82170 9414 82226
rect 9482 82170 9538 82226
rect 9606 82170 9662 82226
rect 9234 82046 9290 82102
rect 9358 82046 9414 82102
rect 9482 82046 9538 82102
rect 9606 82046 9662 82102
rect 9234 81922 9290 81978
rect 9358 81922 9414 81978
rect 9482 81922 9538 81978
rect 9606 81922 9662 81978
rect 9234 64294 9290 64350
rect 9358 64294 9414 64350
rect 9482 64294 9538 64350
rect 9606 64294 9662 64350
rect 9234 64170 9290 64226
rect 9358 64170 9414 64226
rect 9482 64170 9538 64226
rect 9606 64170 9662 64226
rect 9234 64046 9290 64102
rect 9358 64046 9414 64102
rect 9482 64046 9538 64102
rect 9606 64046 9662 64102
rect 9234 63922 9290 63978
rect 9358 63922 9414 63978
rect 9482 63922 9538 63978
rect 9606 63922 9662 63978
rect 9234 46294 9290 46350
rect 9358 46294 9414 46350
rect 9482 46294 9538 46350
rect 9606 46294 9662 46350
rect 9234 46170 9290 46226
rect 9358 46170 9414 46226
rect 9482 46170 9538 46226
rect 9606 46170 9662 46226
rect 9234 46046 9290 46102
rect 9358 46046 9414 46102
rect 9482 46046 9538 46102
rect 9606 46046 9662 46102
rect 9234 45922 9290 45978
rect 9358 45922 9414 45978
rect 9482 45922 9538 45978
rect 9606 45922 9662 45978
rect 9234 28294 9290 28350
rect 9358 28294 9414 28350
rect 9482 28294 9538 28350
rect 9606 28294 9662 28350
rect 9234 28170 9290 28226
rect 9358 28170 9414 28226
rect 9482 28170 9538 28226
rect 9606 28170 9662 28226
rect 9234 28046 9290 28102
rect 9358 28046 9414 28102
rect 9482 28046 9538 28102
rect 9606 28046 9662 28102
rect 9234 27922 9290 27978
rect 9358 27922 9414 27978
rect 9482 27922 9538 27978
rect 9606 27922 9662 27978
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 597156 36290 597212
rect 36358 597156 36414 597212
rect 36482 597156 36538 597212
rect 36606 597156 36662 597212
rect 36234 597032 36290 597088
rect 36358 597032 36414 597088
rect 36482 597032 36538 597088
rect 36606 597032 36662 597088
rect 36234 596908 36290 596964
rect 36358 596908 36414 596964
rect 36482 596908 36538 596964
rect 36606 596908 36662 596964
rect 36234 596784 36290 596840
rect 36358 596784 36414 596840
rect 36482 596784 36538 596840
rect 36606 596784 36662 596840
rect 36234 580294 36290 580350
rect 36358 580294 36414 580350
rect 36482 580294 36538 580350
rect 36606 580294 36662 580350
rect 36234 580170 36290 580226
rect 36358 580170 36414 580226
rect 36482 580170 36538 580226
rect 36606 580170 36662 580226
rect 36234 580046 36290 580102
rect 36358 580046 36414 580102
rect 36482 580046 36538 580102
rect 36606 580046 36662 580102
rect 36234 579922 36290 579978
rect 36358 579922 36414 579978
rect 36482 579922 36538 579978
rect 36606 579922 36662 579978
rect 36234 562294 36290 562350
rect 36358 562294 36414 562350
rect 36482 562294 36538 562350
rect 36606 562294 36662 562350
rect 36234 562170 36290 562226
rect 36358 562170 36414 562226
rect 36482 562170 36538 562226
rect 36606 562170 36662 562226
rect 36234 562046 36290 562102
rect 36358 562046 36414 562102
rect 36482 562046 36538 562102
rect 36606 562046 36662 562102
rect 36234 561922 36290 561978
rect 36358 561922 36414 561978
rect 36482 561922 36538 561978
rect 36606 561922 36662 561978
rect 36234 544294 36290 544350
rect 36358 544294 36414 544350
rect 36482 544294 36538 544350
rect 36606 544294 36662 544350
rect 36234 544170 36290 544226
rect 36358 544170 36414 544226
rect 36482 544170 36538 544226
rect 36606 544170 36662 544226
rect 36234 544046 36290 544102
rect 36358 544046 36414 544102
rect 36482 544046 36538 544102
rect 36606 544046 36662 544102
rect 36234 543922 36290 543978
rect 36358 543922 36414 543978
rect 36482 543922 36538 543978
rect 36606 543922 36662 543978
rect 36234 526294 36290 526350
rect 36358 526294 36414 526350
rect 36482 526294 36538 526350
rect 36606 526294 36662 526350
rect 36234 526170 36290 526226
rect 36358 526170 36414 526226
rect 36482 526170 36538 526226
rect 36606 526170 36662 526226
rect 36234 526046 36290 526102
rect 36358 526046 36414 526102
rect 36482 526046 36538 526102
rect 36606 526046 36662 526102
rect 36234 525922 36290 525978
rect 36358 525922 36414 525978
rect 36482 525922 36538 525978
rect 36606 525922 36662 525978
rect 36234 508294 36290 508350
rect 36358 508294 36414 508350
rect 36482 508294 36538 508350
rect 36606 508294 36662 508350
rect 36234 508170 36290 508226
rect 36358 508170 36414 508226
rect 36482 508170 36538 508226
rect 36606 508170 36662 508226
rect 36234 508046 36290 508102
rect 36358 508046 36414 508102
rect 36482 508046 36538 508102
rect 36606 508046 36662 508102
rect 36234 507922 36290 507978
rect 36358 507922 36414 507978
rect 36482 507922 36538 507978
rect 36606 507922 36662 507978
rect 36234 490294 36290 490350
rect 36358 490294 36414 490350
rect 36482 490294 36538 490350
rect 36606 490294 36662 490350
rect 36234 490170 36290 490226
rect 36358 490170 36414 490226
rect 36482 490170 36538 490226
rect 36606 490170 36662 490226
rect 36234 490046 36290 490102
rect 36358 490046 36414 490102
rect 36482 490046 36538 490102
rect 36606 490046 36662 490102
rect 36234 489922 36290 489978
rect 36358 489922 36414 489978
rect 36482 489922 36538 489978
rect 36606 489922 36662 489978
rect 36234 472294 36290 472350
rect 36358 472294 36414 472350
rect 36482 472294 36538 472350
rect 36606 472294 36662 472350
rect 36234 472170 36290 472226
rect 36358 472170 36414 472226
rect 36482 472170 36538 472226
rect 36606 472170 36662 472226
rect 36234 472046 36290 472102
rect 36358 472046 36414 472102
rect 36482 472046 36538 472102
rect 36606 472046 36662 472102
rect 36234 471922 36290 471978
rect 36358 471922 36414 471978
rect 36482 471922 36538 471978
rect 36606 471922 36662 471978
rect 36234 454294 36290 454350
rect 36358 454294 36414 454350
rect 36482 454294 36538 454350
rect 36606 454294 36662 454350
rect 36234 454170 36290 454226
rect 36358 454170 36414 454226
rect 36482 454170 36538 454226
rect 36606 454170 36662 454226
rect 36234 454046 36290 454102
rect 36358 454046 36414 454102
rect 36482 454046 36538 454102
rect 36606 454046 36662 454102
rect 36234 453922 36290 453978
rect 36358 453922 36414 453978
rect 36482 453922 36538 453978
rect 36606 453922 36662 453978
rect 36234 436294 36290 436350
rect 36358 436294 36414 436350
rect 36482 436294 36538 436350
rect 36606 436294 36662 436350
rect 36234 436170 36290 436226
rect 36358 436170 36414 436226
rect 36482 436170 36538 436226
rect 36606 436170 36662 436226
rect 36234 436046 36290 436102
rect 36358 436046 36414 436102
rect 36482 436046 36538 436102
rect 36606 436046 36662 436102
rect 36234 435922 36290 435978
rect 36358 435922 36414 435978
rect 36482 435922 36538 435978
rect 36606 435922 36662 435978
rect 36234 418294 36290 418350
rect 36358 418294 36414 418350
rect 36482 418294 36538 418350
rect 36606 418294 36662 418350
rect 36234 418170 36290 418226
rect 36358 418170 36414 418226
rect 36482 418170 36538 418226
rect 36606 418170 36662 418226
rect 36234 418046 36290 418102
rect 36358 418046 36414 418102
rect 36482 418046 36538 418102
rect 36606 418046 36662 418102
rect 36234 417922 36290 417978
rect 36358 417922 36414 417978
rect 36482 417922 36538 417978
rect 36606 417922 36662 417978
rect 36234 400294 36290 400350
rect 36358 400294 36414 400350
rect 36482 400294 36538 400350
rect 36606 400294 36662 400350
rect 36234 400170 36290 400226
rect 36358 400170 36414 400226
rect 36482 400170 36538 400226
rect 36606 400170 36662 400226
rect 36234 400046 36290 400102
rect 36358 400046 36414 400102
rect 36482 400046 36538 400102
rect 36606 400046 36662 400102
rect 36234 399922 36290 399978
rect 36358 399922 36414 399978
rect 36482 399922 36538 399978
rect 36606 399922 36662 399978
rect 36234 382294 36290 382350
rect 36358 382294 36414 382350
rect 36482 382294 36538 382350
rect 36606 382294 36662 382350
rect 36234 382170 36290 382226
rect 36358 382170 36414 382226
rect 36482 382170 36538 382226
rect 36606 382170 36662 382226
rect 36234 382046 36290 382102
rect 36358 382046 36414 382102
rect 36482 382046 36538 382102
rect 36606 382046 36662 382102
rect 36234 381922 36290 381978
rect 36358 381922 36414 381978
rect 36482 381922 36538 381978
rect 36606 381922 36662 381978
rect 36234 364294 36290 364350
rect 36358 364294 36414 364350
rect 36482 364294 36538 364350
rect 36606 364294 36662 364350
rect 36234 364170 36290 364226
rect 36358 364170 36414 364226
rect 36482 364170 36538 364226
rect 36606 364170 36662 364226
rect 36234 364046 36290 364102
rect 36358 364046 36414 364102
rect 36482 364046 36538 364102
rect 36606 364046 36662 364102
rect 36234 363922 36290 363978
rect 36358 363922 36414 363978
rect 36482 363922 36538 363978
rect 36606 363922 36662 363978
rect 36234 346294 36290 346350
rect 36358 346294 36414 346350
rect 36482 346294 36538 346350
rect 36606 346294 36662 346350
rect 36234 346170 36290 346226
rect 36358 346170 36414 346226
rect 36482 346170 36538 346226
rect 36606 346170 36662 346226
rect 36234 346046 36290 346102
rect 36358 346046 36414 346102
rect 36482 346046 36538 346102
rect 36606 346046 36662 346102
rect 36234 345922 36290 345978
rect 36358 345922 36414 345978
rect 36482 345922 36538 345978
rect 36606 345922 36662 345978
rect 36234 328294 36290 328350
rect 36358 328294 36414 328350
rect 36482 328294 36538 328350
rect 36606 328294 36662 328350
rect 36234 328170 36290 328226
rect 36358 328170 36414 328226
rect 36482 328170 36538 328226
rect 36606 328170 36662 328226
rect 36234 328046 36290 328102
rect 36358 328046 36414 328102
rect 36482 328046 36538 328102
rect 36606 328046 36662 328102
rect 36234 327922 36290 327978
rect 36358 327922 36414 327978
rect 36482 327922 36538 327978
rect 36606 327922 36662 327978
rect 36234 310294 36290 310350
rect 36358 310294 36414 310350
rect 36482 310294 36538 310350
rect 36606 310294 36662 310350
rect 36234 310170 36290 310226
rect 36358 310170 36414 310226
rect 36482 310170 36538 310226
rect 36606 310170 36662 310226
rect 36234 310046 36290 310102
rect 36358 310046 36414 310102
rect 36482 310046 36538 310102
rect 36606 310046 36662 310102
rect 36234 309922 36290 309978
rect 36358 309922 36414 309978
rect 36482 309922 36538 309978
rect 36606 309922 36662 309978
rect 36234 292294 36290 292350
rect 36358 292294 36414 292350
rect 36482 292294 36538 292350
rect 36606 292294 36662 292350
rect 36234 292170 36290 292226
rect 36358 292170 36414 292226
rect 36482 292170 36538 292226
rect 36606 292170 36662 292226
rect 36234 292046 36290 292102
rect 36358 292046 36414 292102
rect 36482 292046 36538 292102
rect 36606 292046 36662 292102
rect 36234 291922 36290 291978
rect 36358 291922 36414 291978
rect 36482 291922 36538 291978
rect 36606 291922 36662 291978
rect 36234 274294 36290 274350
rect 36358 274294 36414 274350
rect 36482 274294 36538 274350
rect 36606 274294 36662 274350
rect 36234 274170 36290 274226
rect 36358 274170 36414 274226
rect 36482 274170 36538 274226
rect 36606 274170 36662 274226
rect 36234 274046 36290 274102
rect 36358 274046 36414 274102
rect 36482 274046 36538 274102
rect 36606 274046 36662 274102
rect 36234 273922 36290 273978
rect 36358 273922 36414 273978
rect 36482 273922 36538 273978
rect 36606 273922 36662 273978
rect 36234 256294 36290 256350
rect 36358 256294 36414 256350
rect 36482 256294 36538 256350
rect 36606 256294 36662 256350
rect 36234 256170 36290 256226
rect 36358 256170 36414 256226
rect 36482 256170 36538 256226
rect 36606 256170 36662 256226
rect 36234 256046 36290 256102
rect 36358 256046 36414 256102
rect 36482 256046 36538 256102
rect 36606 256046 36662 256102
rect 36234 255922 36290 255978
rect 36358 255922 36414 255978
rect 36482 255922 36538 255978
rect 36606 255922 36662 255978
rect 36234 238294 36290 238350
rect 36358 238294 36414 238350
rect 36482 238294 36538 238350
rect 36606 238294 36662 238350
rect 36234 238170 36290 238226
rect 36358 238170 36414 238226
rect 36482 238170 36538 238226
rect 36606 238170 36662 238226
rect 36234 238046 36290 238102
rect 36358 238046 36414 238102
rect 36482 238046 36538 238102
rect 36606 238046 36662 238102
rect 36234 237922 36290 237978
rect 36358 237922 36414 237978
rect 36482 237922 36538 237978
rect 36606 237922 36662 237978
rect 36234 220294 36290 220350
rect 36358 220294 36414 220350
rect 36482 220294 36538 220350
rect 36606 220294 36662 220350
rect 36234 220170 36290 220226
rect 36358 220170 36414 220226
rect 36482 220170 36538 220226
rect 36606 220170 36662 220226
rect 36234 220046 36290 220102
rect 36358 220046 36414 220102
rect 36482 220046 36538 220102
rect 36606 220046 36662 220102
rect 36234 219922 36290 219978
rect 36358 219922 36414 219978
rect 36482 219922 36538 219978
rect 36606 219922 36662 219978
rect 36234 202294 36290 202350
rect 36358 202294 36414 202350
rect 36482 202294 36538 202350
rect 36606 202294 36662 202350
rect 36234 202170 36290 202226
rect 36358 202170 36414 202226
rect 36482 202170 36538 202226
rect 36606 202170 36662 202226
rect 36234 202046 36290 202102
rect 36358 202046 36414 202102
rect 36482 202046 36538 202102
rect 36606 202046 36662 202102
rect 36234 201922 36290 201978
rect 36358 201922 36414 201978
rect 36482 201922 36538 201978
rect 36606 201922 36662 201978
rect 36234 184294 36290 184350
rect 36358 184294 36414 184350
rect 36482 184294 36538 184350
rect 36606 184294 36662 184350
rect 36234 184170 36290 184226
rect 36358 184170 36414 184226
rect 36482 184170 36538 184226
rect 36606 184170 36662 184226
rect 36234 184046 36290 184102
rect 36358 184046 36414 184102
rect 36482 184046 36538 184102
rect 36606 184046 36662 184102
rect 36234 183922 36290 183978
rect 36358 183922 36414 183978
rect 36482 183922 36538 183978
rect 36606 183922 36662 183978
rect 36234 166294 36290 166350
rect 36358 166294 36414 166350
rect 36482 166294 36538 166350
rect 36606 166294 36662 166350
rect 36234 166170 36290 166226
rect 36358 166170 36414 166226
rect 36482 166170 36538 166226
rect 36606 166170 36662 166226
rect 36234 166046 36290 166102
rect 36358 166046 36414 166102
rect 36482 166046 36538 166102
rect 36606 166046 36662 166102
rect 36234 165922 36290 165978
rect 36358 165922 36414 165978
rect 36482 165922 36538 165978
rect 36606 165922 36662 165978
rect 36234 148294 36290 148350
rect 36358 148294 36414 148350
rect 36482 148294 36538 148350
rect 36606 148294 36662 148350
rect 36234 148170 36290 148226
rect 36358 148170 36414 148226
rect 36482 148170 36538 148226
rect 36606 148170 36662 148226
rect 36234 148046 36290 148102
rect 36358 148046 36414 148102
rect 36482 148046 36538 148102
rect 36606 148046 36662 148102
rect 36234 147922 36290 147978
rect 36358 147922 36414 147978
rect 36482 147922 36538 147978
rect 36606 147922 36662 147978
rect 36234 130294 36290 130350
rect 36358 130294 36414 130350
rect 36482 130294 36538 130350
rect 36606 130294 36662 130350
rect 36234 130170 36290 130226
rect 36358 130170 36414 130226
rect 36482 130170 36538 130226
rect 36606 130170 36662 130226
rect 36234 130046 36290 130102
rect 36358 130046 36414 130102
rect 36482 130046 36538 130102
rect 36606 130046 36662 130102
rect 36234 129922 36290 129978
rect 36358 129922 36414 129978
rect 36482 129922 36538 129978
rect 36606 129922 36662 129978
rect 36234 112294 36290 112350
rect 36358 112294 36414 112350
rect 36482 112294 36538 112350
rect 36606 112294 36662 112350
rect 36234 112170 36290 112226
rect 36358 112170 36414 112226
rect 36482 112170 36538 112226
rect 36606 112170 36662 112226
rect 36234 112046 36290 112102
rect 36358 112046 36414 112102
rect 36482 112046 36538 112102
rect 36606 112046 36662 112102
rect 36234 111922 36290 111978
rect 36358 111922 36414 111978
rect 36482 111922 36538 111978
rect 36606 111922 36662 111978
rect 36234 94294 36290 94350
rect 36358 94294 36414 94350
rect 36482 94294 36538 94350
rect 36606 94294 36662 94350
rect 36234 94170 36290 94226
rect 36358 94170 36414 94226
rect 36482 94170 36538 94226
rect 36606 94170 36662 94226
rect 36234 94046 36290 94102
rect 36358 94046 36414 94102
rect 36482 94046 36538 94102
rect 36606 94046 36662 94102
rect 36234 93922 36290 93978
rect 36358 93922 36414 93978
rect 36482 93922 36538 93978
rect 36606 93922 36662 93978
rect 36234 76294 36290 76350
rect 36358 76294 36414 76350
rect 36482 76294 36538 76350
rect 36606 76294 36662 76350
rect 36234 76170 36290 76226
rect 36358 76170 36414 76226
rect 36482 76170 36538 76226
rect 36606 76170 36662 76226
rect 36234 76046 36290 76102
rect 36358 76046 36414 76102
rect 36482 76046 36538 76102
rect 36606 76046 36662 76102
rect 36234 75922 36290 75978
rect 36358 75922 36414 75978
rect 36482 75922 36538 75978
rect 36606 75922 36662 75978
rect 36234 58294 36290 58350
rect 36358 58294 36414 58350
rect 36482 58294 36538 58350
rect 36606 58294 36662 58350
rect 36234 58170 36290 58226
rect 36358 58170 36414 58226
rect 36482 58170 36538 58226
rect 36606 58170 36662 58226
rect 36234 58046 36290 58102
rect 36358 58046 36414 58102
rect 36482 58046 36538 58102
rect 36606 58046 36662 58102
rect 36234 57922 36290 57978
rect 36358 57922 36414 57978
rect 36482 57922 36538 57978
rect 36606 57922 36662 57978
rect 36234 40294 36290 40350
rect 36358 40294 36414 40350
rect 36482 40294 36538 40350
rect 36606 40294 36662 40350
rect 36234 40170 36290 40226
rect 36358 40170 36414 40226
rect 36482 40170 36538 40226
rect 36606 40170 36662 40226
rect 36234 40046 36290 40102
rect 36358 40046 36414 40102
rect 36482 40046 36538 40102
rect 36606 40046 36662 40102
rect 36234 39922 36290 39978
rect 36358 39922 36414 39978
rect 36482 39922 36538 39978
rect 36606 39922 36662 39978
rect 36234 22294 36290 22350
rect 36358 22294 36414 22350
rect 36482 22294 36538 22350
rect 36606 22294 36662 22350
rect 36234 22170 36290 22226
rect 36358 22170 36414 22226
rect 36482 22170 36538 22226
rect 36606 22170 36662 22226
rect 36234 22046 36290 22102
rect 36358 22046 36414 22102
rect 36482 22046 36538 22102
rect 36606 22046 36662 22102
rect 36234 21922 36290 21978
rect 36358 21922 36414 21978
rect 36482 21922 36538 21978
rect 36606 21922 36662 21978
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 66954 597156 67010 597212
rect 67078 597156 67134 597212
rect 67202 597156 67258 597212
rect 67326 597156 67382 597212
rect 66954 597032 67010 597088
rect 67078 597032 67134 597088
rect 67202 597032 67258 597088
rect 67326 597032 67382 597088
rect 66954 596908 67010 596964
rect 67078 596908 67134 596964
rect 67202 596908 67258 596964
rect 67326 596908 67382 596964
rect 66954 596784 67010 596840
rect 67078 596784 67134 596840
rect 67202 596784 67258 596840
rect 67326 596784 67382 596840
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 39954 568294 40010 568350
rect 40078 568294 40134 568350
rect 40202 568294 40258 568350
rect 40326 568294 40382 568350
rect 39954 568170 40010 568226
rect 40078 568170 40134 568226
rect 40202 568170 40258 568226
rect 40326 568170 40382 568226
rect 39954 568046 40010 568102
rect 40078 568046 40134 568102
rect 40202 568046 40258 568102
rect 40326 568046 40382 568102
rect 39954 567922 40010 567978
rect 40078 567922 40134 567978
rect 40202 567922 40258 567978
rect 40326 567922 40382 567978
rect 39954 550294 40010 550350
rect 40078 550294 40134 550350
rect 40202 550294 40258 550350
rect 40326 550294 40382 550350
rect 39954 550170 40010 550226
rect 40078 550170 40134 550226
rect 40202 550170 40258 550226
rect 40326 550170 40382 550226
rect 39954 550046 40010 550102
rect 40078 550046 40134 550102
rect 40202 550046 40258 550102
rect 40326 550046 40382 550102
rect 39954 549922 40010 549978
rect 40078 549922 40134 549978
rect 40202 549922 40258 549978
rect 40326 549922 40382 549978
rect 39954 532294 40010 532350
rect 40078 532294 40134 532350
rect 40202 532294 40258 532350
rect 40326 532294 40382 532350
rect 39954 532170 40010 532226
rect 40078 532170 40134 532226
rect 40202 532170 40258 532226
rect 40326 532170 40382 532226
rect 39954 532046 40010 532102
rect 40078 532046 40134 532102
rect 40202 532046 40258 532102
rect 40326 532046 40382 532102
rect 39954 531922 40010 531978
rect 40078 531922 40134 531978
rect 40202 531922 40258 531978
rect 40326 531922 40382 531978
rect 39954 514294 40010 514350
rect 40078 514294 40134 514350
rect 40202 514294 40258 514350
rect 40326 514294 40382 514350
rect 39954 514170 40010 514226
rect 40078 514170 40134 514226
rect 40202 514170 40258 514226
rect 40326 514170 40382 514226
rect 39954 514046 40010 514102
rect 40078 514046 40134 514102
rect 40202 514046 40258 514102
rect 40326 514046 40382 514102
rect 39954 513922 40010 513978
rect 40078 513922 40134 513978
rect 40202 513922 40258 513978
rect 40326 513922 40382 513978
rect 39954 496294 40010 496350
rect 40078 496294 40134 496350
rect 40202 496294 40258 496350
rect 40326 496294 40382 496350
rect 39954 496170 40010 496226
rect 40078 496170 40134 496226
rect 40202 496170 40258 496226
rect 40326 496170 40382 496226
rect 39954 496046 40010 496102
rect 40078 496046 40134 496102
rect 40202 496046 40258 496102
rect 40326 496046 40382 496102
rect 39954 495922 40010 495978
rect 40078 495922 40134 495978
rect 40202 495922 40258 495978
rect 40326 495922 40382 495978
rect 39954 478294 40010 478350
rect 40078 478294 40134 478350
rect 40202 478294 40258 478350
rect 40326 478294 40382 478350
rect 39954 478170 40010 478226
rect 40078 478170 40134 478226
rect 40202 478170 40258 478226
rect 40326 478170 40382 478226
rect 39954 478046 40010 478102
rect 40078 478046 40134 478102
rect 40202 478046 40258 478102
rect 40326 478046 40382 478102
rect 39954 477922 40010 477978
rect 40078 477922 40134 477978
rect 40202 477922 40258 477978
rect 40326 477922 40382 477978
rect 39954 460294 40010 460350
rect 40078 460294 40134 460350
rect 40202 460294 40258 460350
rect 40326 460294 40382 460350
rect 39954 460170 40010 460226
rect 40078 460170 40134 460226
rect 40202 460170 40258 460226
rect 40326 460170 40382 460226
rect 39954 460046 40010 460102
rect 40078 460046 40134 460102
rect 40202 460046 40258 460102
rect 40326 460046 40382 460102
rect 39954 459922 40010 459978
rect 40078 459922 40134 459978
rect 40202 459922 40258 459978
rect 40326 459922 40382 459978
rect 39954 442294 40010 442350
rect 40078 442294 40134 442350
rect 40202 442294 40258 442350
rect 40326 442294 40382 442350
rect 39954 442170 40010 442226
rect 40078 442170 40134 442226
rect 40202 442170 40258 442226
rect 40326 442170 40382 442226
rect 39954 442046 40010 442102
rect 40078 442046 40134 442102
rect 40202 442046 40258 442102
rect 40326 442046 40382 442102
rect 39954 441922 40010 441978
rect 40078 441922 40134 441978
rect 40202 441922 40258 441978
rect 40326 441922 40382 441978
rect 39954 424294 40010 424350
rect 40078 424294 40134 424350
rect 40202 424294 40258 424350
rect 40326 424294 40382 424350
rect 39954 424170 40010 424226
rect 40078 424170 40134 424226
rect 40202 424170 40258 424226
rect 40326 424170 40382 424226
rect 39954 424046 40010 424102
rect 40078 424046 40134 424102
rect 40202 424046 40258 424102
rect 40326 424046 40382 424102
rect 39954 423922 40010 423978
rect 40078 423922 40134 423978
rect 40202 423922 40258 423978
rect 40326 423922 40382 423978
rect 39954 406294 40010 406350
rect 40078 406294 40134 406350
rect 40202 406294 40258 406350
rect 40326 406294 40382 406350
rect 39954 406170 40010 406226
rect 40078 406170 40134 406226
rect 40202 406170 40258 406226
rect 40326 406170 40382 406226
rect 39954 406046 40010 406102
rect 40078 406046 40134 406102
rect 40202 406046 40258 406102
rect 40326 406046 40382 406102
rect 39954 405922 40010 405978
rect 40078 405922 40134 405978
rect 40202 405922 40258 405978
rect 40326 405922 40382 405978
rect 39954 388294 40010 388350
rect 40078 388294 40134 388350
rect 40202 388294 40258 388350
rect 40326 388294 40382 388350
rect 39954 388170 40010 388226
rect 40078 388170 40134 388226
rect 40202 388170 40258 388226
rect 40326 388170 40382 388226
rect 39954 388046 40010 388102
rect 40078 388046 40134 388102
rect 40202 388046 40258 388102
rect 40326 388046 40382 388102
rect 39954 387922 40010 387978
rect 40078 387922 40134 387978
rect 40202 387922 40258 387978
rect 40326 387922 40382 387978
rect 39954 370294 40010 370350
rect 40078 370294 40134 370350
rect 40202 370294 40258 370350
rect 40326 370294 40382 370350
rect 39954 370170 40010 370226
rect 40078 370170 40134 370226
rect 40202 370170 40258 370226
rect 40326 370170 40382 370226
rect 39954 370046 40010 370102
rect 40078 370046 40134 370102
rect 40202 370046 40258 370102
rect 40326 370046 40382 370102
rect 39954 369922 40010 369978
rect 40078 369922 40134 369978
rect 40202 369922 40258 369978
rect 40326 369922 40382 369978
rect 39954 352294 40010 352350
rect 40078 352294 40134 352350
rect 40202 352294 40258 352350
rect 40326 352294 40382 352350
rect 39954 352170 40010 352226
rect 40078 352170 40134 352226
rect 40202 352170 40258 352226
rect 40326 352170 40382 352226
rect 39954 352046 40010 352102
rect 40078 352046 40134 352102
rect 40202 352046 40258 352102
rect 40326 352046 40382 352102
rect 39954 351922 40010 351978
rect 40078 351922 40134 351978
rect 40202 351922 40258 351978
rect 40326 351922 40382 351978
rect 39954 334294 40010 334350
rect 40078 334294 40134 334350
rect 40202 334294 40258 334350
rect 40326 334294 40382 334350
rect 39954 334170 40010 334226
rect 40078 334170 40134 334226
rect 40202 334170 40258 334226
rect 40326 334170 40382 334226
rect 39954 334046 40010 334102
rect 40078 334046 40134 334102
rect 40202 334046 40258 334102
rect 40326 334046 40382 334102
rect 39954 333922 40010 333978
rect 40078 333922 40134 333978
rect 40202 333922 40258 333978
rect 40326 333922 40382 333978
rect 39954 316294 40010 316350
rect 40078 316294 40134 316350
rect 40202 316294 40258 316350
rect 40326 316294 40382 316350
rect 39954 316170 40010 316226
rect 40078 316170 40134 316226
rect 40202 316170 40258 316226
rect 40326 316170 40382 316226
rect 39954 316046 40010 316102
rect 40078 316046 40134 316102
rect 40202 316046 40258 316102
rect 40326 316046 40382 316102
rect 39954 315922 40010 315978
rect 40078 315922 40134 315978
rect 40202 315922 40258 315978
rect 40326 315922 40382 315978
rect 66954 580294 67010 580350
rect 67078 580294 67134 580350
rect 67202 580294 67258 580350
rect 67326 580294 67382 580350
rect 66954 580170 67010 580226
rect 67078 580170 67134 580226
rect 67202 580170 67258 580226
rect 67326 580170 67382 580226
rect 66954 580046 67010 580102
rect 67078 580046 67134 580102
rect 67202 580046 67258 580102
rect 67326 580046 67382 580102
rect 66954 579922 67010 579978
rect 67078 579922 67134 579978
rect 67202 579922 67258 579978
rect 67326 579922 67382 579978
rect 66954 562294 67010 562350
rect 67078 562294 67134 562350
rect 67202 562294 67258 562350
rect 67326 562294 67382 562350
rect 66954 562170 67010 562226
rect 67078 562170 67134 562226
rect 67202 562170 67258 562226
rect 67326 562170 67382 562226
rect 66954 562046 67010 562102
rect 67078 562046 67134 562102
rect 67202 562046 67258 562102
rect 67326 562046 67382 562102
rect 66954 561922 67010 561978
rect 67078 561922 67134 561978
rect 67202 561922 67258 561978
rect 67326 561922 67382 561978
rect 55356 551042 55412 551098
rect 53116 300662 53172 300718
rect 39954 298294 40010 298350
rect 40078 298294 40134 298350
rect 40202 298294 40258 298350
rect 40326 298294 40382 298350
rect 39954 298170 40010 298226
rect 40078 298170 40134 298226
rect 40202 298170 40258 298226
rect 40326 298170 40382 298226
rect 39954 298046 40010 298102
rect 40078 298046 40134 298102
rect 40202 298046 40258 298102
rect 40326 298046 40382 298102
rect 39954 297922 40010 297978
rect 40078 297922 40134 297978
rect 40202 297922 40258 297978
rect 40326 297922 40382 297978
rect 53228 293642 53284 293698
rect 53564 296882 53620 296938
rect 54348 300302 54404 300358
rect 53676 291662 53732 291718
rect 54572 288422 54628 288478
rect 53452 287162 53508 287218
rect 53340 285362 53396 285418
rect 54796 290582 54852 290638
rect 55020 290222 55076 290278
rect 55132 282122 55188 282178
rect 39954 280294 40010 280350
rect 40078 280294 40134 280350
rect 40202 280294 40258 280350
rect 40326 280294 40382 280350
rect 39954 280170 40010 280226
rect 40078 280170 40134 280226
rect 40202 280170 40258 280226
rect 40326 280170 40382 280226
rect 39954 280046 40010 280102
rect 40078 280046 40134 280102
rect 40202 280046 40258 280102
rect 40326 280046 40382 280102
rect 39954 279922 40010 279978
rect 40078 279922 40134 279978
rect 40202 279922 40258 279978
rect 40326 279922 40382 279978
rect 39954 262294 40010 262350
rect 40078 262294 40134 262350
rect 40202 262294 40258 262350
rect 40326 262294 40382 262350
rect 39954 262170 40010 262226
rect 40078 262170 40134 262226
rect 40202 262170 40258 262226
rect 40326 262170 40382 262226
rect 39954 262046 40010 262102
rect 40078 262046 40134 262102
rect 40202 262046 40258 262102
rect 40326 262046 40382 262102
rect 39954 261922 40010 261978
rect 40078 261922 40134 261978
rect 40202 261922 40258 261978
rect 40326 261922 40382 261978
rect 39954 244294 40010 244350
rect 40078 244294 40134 244350
rect 40202 244294 40258 244350
rect 40326 244294 40382 244350
rect 39954 244170 40010 244226
rect 40078 244170 40134 244226
rect 40202 244170 40258 244226
rect 40326 244170 40382 244226
rect 39954 244046 40010 244102
rect 40078 244046 40134 244102
rect 40202 244046 40258 244102
rect 40326 244046 40382 244102
rect 39954 243922 40010 243978
rect 40078 243922 40134 243978
rect 40202 243922 40258 243978
rect 40326 243922 40382 243978
rect 39954 226294 40010 226350
rect 40078 226294 40134 226350
rect 40202 226294 40258 226350
rect 40326 226294 40382 226350
rect 39954 226170 40010 226226
rect 40078 226170 40134 226226
rect 40202 226170 40258 226226
rect 40326 226170 40382 226226
rect 39954 226046 40010 226102
rect 40078 226046 40134 226102
rect 40202 226046 40258 226102
rect 40326 226046 40382 226102
rect 39954 225922 40010 225978
rect 40078 225922 40134 225978
rect 40202 225922 40258 225978
rect 40326 225922 40382 225978
rect 39954 208294 40010 208350
rect 40078 208294 40134 208350
rect 40202 208294 40258 208350
rect 40326 208294 40382 208350
rect 39954 208170 40010 208226
rect 40078 208170 40134 208226
rect 40202 208170 40258 208226
rect 40326 208170 40382 208226
rect 39954 208046 40010 208102
rect 40078 208046 40134 208102
rect 40202 208046 40258 208102
rect 40326 208046 40382 208102
rect 39954 207922 40010 207978
rect 40078 207922 40134 207978
rect 40202 207922 40258 207978
rect 40326 207922 40382 207978
rect 39954 190294 40010 190350
rect 40078 190294 40134 190350
rect 40202 190294 40258 190350
rect 40326 190294 40382 190350
rect 39954 190170 40010 190226
rect 40078 190170 40134 190226
rect 40202 190170 40258 190226
rect 40326 190170 40382 190226
rect 39954 190046 40010 190102
rect 40078 190046 40134 190102
rect 40202 190046 40258 190102
rect 40326 190046 40382 190102
rect 39954 189922 40010 189978
rect 40078 189922 40134 189978
rect 40202 189922 40258 189978
rect 40326 189922 40382 189978
rect 39954 172294 40010 172350
rect 40078 172294 40134 172350
rect 40202 172294 40258 172350
rect 40326 172294 40382 172350
rect 39954 172170 40010 172226
rect 40078 172170 40134 172226
rect 40202 172170 40258 172226
rect 40326 172170 40382 172226
rect 39954 172046 40010 172102
rect 40078 172046 40134 172102
rect 40202 172046 40258 172102
rect 40326 172046 40382 172102
rect 39954 171922 40010 171978
rect 40078 171922 40134 171978
rect 40202 171922 40258 171978
rect 40326 171922 40382 171978
rect 39954 154294 40010 154350
rect 40078 154294 40134 154350
rect 40202 154294 40258 154350
rect 40326 154294 40382 154350
rect 39954 154170 40010 154226
rect 40078 154170 40134 154226
rect 40202 154170 40258 154226
rect 40326 154170 40382 154226
rect 39954 154046 40010 154102
rect 40078 154046 40134 154102
rect 40202 154046 40258 154102
rect 40326 154046 40382 154102
rect 39954 153922 40010 153978
rect 40078 153922 40134 153978
rect 40202 153922 40258 153978
rect 40326 153922 40382 153978
rect 58716 547802 58772 547858
rect 56588 427202 56644 427258
rect 57036 427022 57092 427078
rect 56700 425042 56756 425098
rect 56812 423422 56868 423478
rect 66954 544294 67010 544350
rect 67078 544294 67134 544350
rect 67202 544294 67258 544350
rect 67326 544294 67382 544350
rect 66954 544170 67010 544226
rect 67078 544170 67134 544226
rect 67202 544170 67258 544226
rect 67326 544170 67382 544226
rect 66954 544046 67010 544102
rect 67078 544046 67134 544102
rect 67202 544046 67258 544102
rect 67326 544046 67382 544102
rect 66954 543922 67010 543978
rect 67078 543922 67134 543978
rect 67202 543922 67258 543978
rect 67326 543922 67382 543978
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 70674 568294 70730 568350
rect 70798 568294 70854 568350
rect 70922 568294 70978 568350
rect 71046 568294 71102 568350
rect 70674 568170 70730 568226
rect 70798 568170 70854 568226
rect 70922 568170 70978 568226
rect 71046 568170 71102 568226
rect 70674 568046 70730 568102
rect 70798 568046 70854 568102
rect 70922 568046 70978 568102
rect 71046 568046 71102 568102
rect 70674 567922 70730 567978
rect 70798 567922 70854 567978
rect 70922 567922 70978 567978
rect 71046 567922 71102 567978
rect 97674 597156 97730 597212
rect 97798 597156 97854 597212
rect 97922 597156 97978 597212
rect 98046 597156 98102 597212
rect 97674 597032 97730 597088
rect 97798 597032 97854 597088
rect 97922 597032 97978 597088
rect 98046 597032 98102 597088
rect 97674 596908 97730 596964
rect 97798 596908 97854 596964
rect 97922 596908 97978 596964
rect 98046 596908 98102 596964
rect 97674 596784 97730 596840
rect 97798 596784 97854 596840
rect 97922 596784 97978 596840
rect 98046 596784 98102 596840
rect 97674 580294 97730 580350
rect 97798 580294 97854 580350
rect 97922 580294 97978 580350
rect 98046 580294 98102 580350
rect 97674 580170 97730 580226
rect 97798 580170 97854 580226
rect 97922 580170 97978 580226
rect 98046 580170 98102 580226
rect 97674 580046 97730 580102
rect 97798 580046 97854 580102
rect 97922 580046 97978 580102
rect 98046 580046 98102 580102
rect 97674 579922 97730 579978
rect 97798 579922 97854 579978
rect 97922 579922 97978 579978
rect 98046 579922 98102 579978
rect 97674 562294 97730 562350
rect 97798 562294 97854 562350
rect 97922 562294 97978 562350
rect 98046 562294 98102 562350
rect 97674 562170 97730 562226
rect 97798 562170 97854 562226
rect 97922 562170 97978 562226
rect 98046 562170 98102 562226
rect 97674 562046 97730 562102
rect 97798 562046 97854 562102
rect 97922 562046 97978 562102
rect 98046 562046 98102 562102
rect 97674 561922 97730 561978
rect 97798 561922 97854 561978
rect 97922 561922 97978 561978
rect 98046 561922 98102 561978
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 101394 568294 101450 568350
rect 101518 568294 101574 568350
rect 101642 568294 101698 568350
rect 101766 568294 101822 568350
rect 101394 568170 101450 568226
rect 101518 568170 101574 568226
rect 101642 568170 101698 568226
rect 101766 568170 101822 568226
rect 101394 568046 101450 568102
rect 101518 568046 101574 568102
rect 101642 568046 101698 568102
rect 101766 568046 101822 568102
rect 101394 567922 101450 567978
rect 101518 567922 101574 567978
rect 101642 567922 101698 567978
rect 101766 567922 101822 567978
rect 128394 597156 128450 597212
rect 128518 597156 128574 597212
rect 128642 597156 128698 597212
rect 128766 597156 128822 597212
rect 128394 597032 128450 597088
rect 128518 597032 128574 597088
rect 128642 597032 128698 597088
rect 128766 597032 128822 597088
rect 128394 596908 128450 596964
rect 128518 596908 128574 596964
rect 128642 596908 128698 596964
rect 128766 596908 128822 596964
rect 128394 596784 128450 596840
rect 128518 596784 128574 596840
rect 128642 596784 128698 596840
rect 128766 596784 128822 596840
rect 128394 580294 128450 580350
rect 128518 580294 128574 580350
rect 128642 580294 128698 580350
rect 128766 580294 128822 580350
rect 128394 580170 128450 580226
rect 128518 580170 128574 580226
rect 128642 580170 128698 580226
rect 128766 580170 128822 580226
rect 128394 580046 128450 580102
rect 128518 580046 128574 580102
rect 128642 580046 128698 580102
rect 128766 580046 128822 580102
rect 128394 579922 128450 579978
rect 128518 579922 128574 579978
rect 128642 579922 128698 579978
rect 128766 579922 128822 579978
rect 128394 562294 128450 562350
rect 128518 562294 128574 562350
rect 128642 562294 128698 562350
rect 128766 562294 128822 562350
rect 128394 562170 128450 562226
rect 128518 562170 128574 562226
rect 128642 562170 128698 562226
rect 128766 562170 128822 562226
rect 128394 562046 128450 562102
rect 128518 562046 128574 562102
rect 128642 562046 128698 562102
rect 128766 562046 128822 562102
rect 128394 561922 128450 561978
rect 128518 561922 128574 561978
rect 128642 561922 128698 561978
rect 128766 561922 128822 561978
rect 70674 550294 70730 550350
rect 70798 550294 70854 550350
rect 70922 550294 70978 550350
rect 71046 550294 71102 550350
rect 70674 550170 70730 550226
rect 70798 550170 70854 550226
rect 70922 550170 70978 550226
rect 71046 550170 71102 550226
rect 70674 550046 70730 550102
rect 70798 550046 70854 550102
rect 70922 550046 70978 550102
rect 71046 550046 71102 550102
rect 70674 549922 70730 549978
rect 70798 549922 70854 549978
rect 70922 549922 70978 549978
rect 71046 549922 71102 549978
rect 121996 547982 122052 548038
rect 94810 544377 94866 544433
rect 94934 544377 94990 544433
rect 94810 544253 94866 544309
rect 94934 544253 94990 544309
rect 95058 544377 95114 544433
rect 95182 544377 95238 544433
rect 95306 544377 95362 544433
rect 95430 544377 95486 544433
rect 95058 544253 95114 544309
rect 95182 544253 95238 544309
rect 95306 544253 95362 544309
rect 95430 544253 95486 544309
rect 95554 544377 95610 544433
rect 95678 544377 95734 544433
rect 95802 544377 95858 544433
rect 95926 544377 95982 544433
rect 95554 544253 95610 544309
rect 95678 544253 95734 544309
rect 95802 544253 95858 544309
rect 95926 544253 95982 544309
rect 96050 544377 96106 544433
rect 96174 544377 96230 544433
rect 96298 544377 96354 544433
rect 96422 544377 96478 544433
rect 96050 544253 96106 544309
rect 96174 544253 96230 544309
rect 96298 544253 96354 544309
rect 96422 544253 96478 544309
rect 96546 544377 96602 544433
rect 96670 544377 96726 544433
rect 96794 544377 96850 544433
rect 96918 544377 96974 544433
rect 96546 544253 96602 544309
rect 96670 544253 96726 544309
rect 96794 544253 96850 544309
rect 96918 544253 96974 544309
rect 97042 544377 97098 544433
rect 97166 544377 97222 544433
rect 97290 544377 97346 544433
rect 97414 544377 97470 544433
rect 97042 544253 97098 544309
rect 97166 544253 97222 544309
rect 97290 544253 97346 544309
rect 97414 544253 97470 544309
rect 97538 544377 97594 544433
rect 97662 544377 97718 544433
rect 97786 544377 97842 544433
rect 97910 544377 97966 544433
rect 97538 544253 97594 544309
rect 97662 544253 97718 544309
rect 97786 544253 97842 544309
rect 97910 544253 97966 544309
rect 98034 544377 98090 544433
rect 98158 544377 98214 544433
rect 98282 544377 98338 544433
rect 98406 544377 98462 544433
rect 98034 544253 98090 544309
rect 98158 544253 98214 544309
rect 98282 544253 98338 544309
rect 98406 544253 98462 544309
rect 98530 544377 98586 544433
rect 98654 544377 98710 544433
rect 98778 544377 98834 544433
rect 98902 544377 98958 544433
rect 98530 544253 98586 544309
rect 98654 544253 98710 544309
rect 98778 544253 98834 544309
rect 98902 544253 98958 544309
rect 99026 544377 99082 544433
rect 99150 544377 99206 544433
rect 99274 544377 99330 544433
rect 99398 544377 99454 544433
rect 99026 544253 99082 544309
rect 99150 544253 99206 544309
rect 99274 544253 99330 544309
rect 99398 544253 99454 544309
rect 99522 544377 99578 544433
rect 99646 544377 99702 544433
rect 99770 544377 99826 544433
rect 99894 544377 99950 544433
rect 99522 544253 99578 544309
rect 99646 544253 99702 544309
rect 99770 544253 99826 544309
rect 99894 544253 99950 544309
rect 100018 544377 100074 544433
rect 100142 544377 100198 544433
rect 100266 544377 100322 544433
rect 100390 544377 100446 544433
rect 100018 544253 100074 544309
rect 100142 544253 100198 544309
rect 100266 544253 100322 544309
rect 100390 544253 100446 544309
rect 100514 544377 100570 544433
rect 100638 544377 100694 544433
rect 100762 544377 100818 544433
rect 100886 544377 100942 544433
rect 100514 544253 100570 544309
rect 100638 544253 100694 544309
rect 100762 544253 100818 544309
rect 100886 544253 100942 544309
rect 101010 544377 101066 544433
rect 101134 544377 101190 544433
rect 101258 544377 101314 544433
rect 101382 544377 101438 544433
rect 101010 544253 101066 544309
rect 101134 544253 101190 544309
rect 101258 544253 101314 544309
rect 101382 544253 101438 544309
rect 101506 544377 101562 544433
rect 101630 544377 101686 544433
rect 101754 544377 101810 544433
rect 101878 544377 101934 544433
rect 101506 544253 101562 544309
rect 101630 544253 101686 544309
rect 101754 544253 101810 544309
rect 101878 544253 101934 544309
rect 102002 544377 102058 544433
rect 102126 544377 102182 544433
rect 102250 544377 102306 544433
rect 102374 544377 102430 544433
rect 102002 544253 102058 544309
rect 102126 544253 102182 544309
rect 102250 544253 102306 544309
rect 102374 544253 102430 544309
rect 102498 544377 102554 544433
rect 102622 544377 102678 544433
rect 102746 544377 102802 544433
rect 102870 544377 102926 544433
rect 102498 544253 102554 544309
rect 102622 544253 102678 544309
rect 102746 544253 102802 544309
rect 102870 544253 102926 544309
rect 102994 544377 103050 544433
rect 103118 544377 103174 544433
rect 103242 544377 103298 544433
rect 103366 544377 103422 544433
rect 102994 544253 103050 544309
rect 103118 544253 103174 544309
rect 103242 544253 103298 544309
rect 103366 544253 103422 544309
rect 103490 544377 103546 544433
rect 103614 544377 103670 544433
rect 103738 544377 103794 544433
rect 103862 544377 103918 544433
rect 103490 544253 103546 544309
rect 103614 544253 103670 544309
rect 103738 544253 103794 544309
rect 103862 544253 103918 544309
rect 103986 544377 104042 544433
rect 104110 544377 104166 544433
rect 104234 544377 104290 544433
rect 104358 544377 104414 544433
rect 103986 544253 104042 544309
rect 104110 544253 104166 544309
rect 104234 544253 104290 544309
rect 104358 544253 104414 544309
rect 104482 544377 104538 544433
rect 104606 544377 104662 544433
rect 104730 544377 104786 544433
rect 104854 544377 104910 544433
rect 104482 544253 104538 544309
rect 104606 544253 104662 544309
rect 104730 544253 104786 544309
rect 104854 544253 104910 544309
rect 104978 544377 105034 544433
rect 105102 544377 105158 544433
rect 105226 544377 105282 544433
rect 105350 544377 105406 544433
rect 104978 544253 105034 544309
rect 105102 544253 105158 544309
rect 105226 544253 105282 544309
rect 105350 544253 105406 544309
rect 105474 544377 105530 544433
rect 105598 544377 105654 544433
rect 105722 544377 105778 544433
rect 105846 544377 105902 544433
rect 105474 544253 105530 544309
rect 105598 544253 105654 544309
rect 105722 544253 105778 544309
rect 105846 544253 105902 544309
rect 105970 544377 106026 544433
rect 106094 544377 106150 544433
rect 106218 544377 106274 544433
rect 106342 544377 106398 544433
rect 105970 544253 106026 544309
rect 106094 544253 106150 544309
rect 106218 544253 106274 544309
rect 106342 544253 106398 544309
rect 106466 544377 106522 544433
rect 106590 544377 106646 544433
rect 106714 544377 106770 544433
rect 106838 544377 106894 544433
rect 106466 544253 106522 544309
rect 106590 544253 106646 544309
rect 106714 544253 106770 544309
rect 106838 544253 106894 544309
rect 106962 544377 107018 544433
rect 107086 544377 107142 544433
rect 107210 544377 107266 544433
rect 107334 544377 107390 544433
rect 106962 544253 107018 544309
rect 107086 544253 107142 544309
rect 107210 544253 107266 544309
rect 107334 544253 107390 544309
rect 94630 544034 94686 544090
rect 94754 544034 94810 544090
rect 94878 544034 94934 544090
rect 95002 544034 95058 544090
rect 95126 544034 95182 544090
rect 95250 544034 95306 544090
rect 95374 544034 95430 544090
rect 95498 544034 95554 544090
rect 95622 544034 95678 544090
rect 95746 544034 95802 544090
rect 95870 544034 95926 544090
rect 95994 544034 96050 544090
rect 96118 544034 96174 544090
rect 96242 544034 96298 544090
rect 96366 544034 96422 544090
rect 96490 544034 96546 544090
rect 96614 544034 96670 544090
rect 96738 544034 96794 544090
rect 96862 544034 96918 544090
rect 96986 544034 97042 544090
rect 97110 544034 97166 544090
rect 97234 544034 97290 544090
rect 97358 544034 97414 544090
rect 97482 544034 97538 544090
rect 97606 544034 97662 544090
rect 97730 544034 97786 544090
rect 97854 544034 97910 544090
rect 97978 544034 98034 544090
rect 98102 544034 98158 544090
rect 98226 544034 98282 544090
rect 98350 544034 98406 544090
rect 98474 544034 98530 544090
rect 98598 544034 98654 544090
rect 98722 544034 98778 544090
rect 98846 544034 98902 544090
rect 98970 544034 99026 544090
rect 99094 544034 99150 544090
rect 99218 544034 99274 544090
rect 99342 544034 99398 544090
rect 99466 544034 99522 544090
rect 99590 544034 99646 544090
rect 99714 544034 99770 544090
rect 99838 544034 99894 544090
rect 99962 544034 100018 544090
rect 100086 544034 100142 544090
rect 100210 544034 100266 544090
rect 100334 544034 100390 544090
rect 100458 544034 100514 544090
rect 100582 544034 100638 544090
rect 100706 544034 100762 544090
rect 100830 544034 100886 544090
rect 100954 544034 101010 544090
rect 101078 544034 101134 544090
rect 101202 544034 101258 544090
rect 101326 544034 101382 544090
rect 101450 544034 101506 544090
rect 101574 544034 101630 544090
rect 101698 544034 101754 544090
rect 101822 544034 101878 544090
rect 101946 544034 102002 544090
rect 102070 544034 102126 544090
rect 102194 544034 102250 544090
rect 102318 544034 102374 544090
rect 102442 544034 102498 544090
rect 102566 544034 102622 544090
rect 102690 544034 102746 544090
rect 102814 544034 102870 544090
rect 102938 544034 102994 544090
rect 103062 544034 103118 544090
rect 103186 544034 103242 544090
rect 103310 544034 103366 544090
rect 103434 544034 103490 544090
rect 103558 544034 103614 544090
rect 103682 544034 103738 544090
rect 103806 544034 103862 544090
rect 103930 544034 103986 544090
rect 104054 544034 104110 544090
rect 104178 544034 104234 544090
rect 104302 544034 104358 544090
rect 104426 544034 104482 544090
rect 104550 544034 104606 544090
rect 104674 544034 104730 544090
rect 104798 544034 104854 544090
rect 104922 544034 104978 544090
rect 105046 544034 105102 544090
rect 105170 544034 105226 544090
rect 105294 544034 105350 544090
rect 105418 544034 105474 544090
rect 105542 544034 105598 544090
rect 105666 544034 105722 544090
rect 105790 544034 105846 544090
rect 105914 544034 105970 544090
rect 106038 544034 106094 544090
rect 106162 544034 106218 544090
rect 106286 544034 106342 544090
rect 106410 544034 106466 544090
rect 106534 544034 106590 544090
rect 106658 544034 106714 544090
rect 106782 544034 106838 544090
rect 106906 544034 106962 544090
rect 107030 544034 107086 544090
rect 107154 544034 107210 544090
rect 94630 543910 94686 543966
rect 94754 543910 94810 543966
rect 94878 543910 94934 543966
rect 95002 543910 95058 543966
rect 95126 543910 95182 543966
rect 95250 543910 95306 543966
rect 95374 543910 95430 543966
rect 95498 543910 95554 543966
rect 95622 543910 95678 543966
rect 95746 543910 95802 543966
rect 95870 543910 95926 543966
rect 95994 543910 96050 543966
rect 96118 543910 96174 543966
rect 96242 543910 96298 543966
rect 96366 543910 96422 543966
rect 96490 543910 96546 543966
rect 96614 543910 96670 543966
rect 96738 543910 96794 543966
rect 96862 543910 96918 543966
rect 96986 543910 97042 543966
rect 97110 543910 97166 543966
rect 97234 543910 97290 543966
rect 97358 543910 97414 543966
rect 97482 543910 97538 543966
rect 97606 543910 97662 543966
rect 97730 543910 97786 543966
rect 97854 543910 97910 543966
rect 97978 543910 98034 543966
rect 98102 543910 98158 543966
rect 98226 543910 98282 543966
rect 98350 543910 98406 543966
rect 98474 543910 98530 543966
rect 98598 543910 98654 543966
rect 98722 543910 98778 543966
rect 98846 543910 98902 543966
rect 98970 543910 99026 543966
rect 99094 543910 99150 543966
rect 99218 543910 99274 543966
rect 99342 543910 99398 543966
rect 99466 543910 99522 543966
rect 99590 543910 99646 543966
rect 99714 543910 99770 543966
rect 99838 543910 99894 543966
rect 99962 543910 100018 543966
rect 100086 543910 100142 543966
rect 100210 543910 100266 543966
rect 100334 543910 100390 543966
rect 100458 543910 100514 543966
rect 100582 543910 100638 543966
rect 100706 543910 100762 543966
rect 100830 543910 100886 543966
rect 100954 543910 101010 543966
rect 101078 543910 101134 543966
rect 101202 543910 101258 543966
rect 101326 543910 101382 543966
rect 101450 543910 101506 543966
rect 101574 543910 101630 543966
rect 101698 543910 101754 543966
rect 101822 543910 101878 543966
rect 101946 543910 102002 543966
rect 102070 543910 102126 543966
rect 102194 543910 102250 543966
rect 102318 543910 102374 543966
rect 102442 543910 102498 543966
rect 102566 543910 102622 543966
rect 102690 543910 102746 543966
rect 102814 543910 102870 543966
rect 102938 543910 102994 543966
rect 103062 543910 103118 543966
rect 103186 543910 103242 543966
rect 103310 543910 103366 543966
rect 103434 543910 103490 543966
rect 103558 543910 103614 543966
rect 103682 543910 103738 543966
rect 103806 543910 103862 543966
rect 103930 543910 103986 543966
rect 104054 543910 104110 543966
rect 104178 543910 104234 543966
rect 104302 543910 104358 543966
rect 104426 543910 104482 543966
rect 104550 543910 104606 543966
rect 104674 543910 104730 543966
rect 104798 543910 104854 543966
rect 104922 543910 104978 543966
rect 105046 543910 105102 543966
rect 105170 543910 105226 543966
rect 105294 543910 105350 543966
rect 105418 543910 105474 543966
rect 105542 543910 105598 543966
rect 105666 543910 105722 543966
rect 105790 543910 105846 543966
rect 105914 543910 105970 543966
rect 106038 543910 106094 543966
rect 106162 543910 106218 543966
rect 106286 543910 106342 543966
rect 106410 543910 106466 543966
rect 106534 543910 106590 543966
rect 106658 543910 106714 543966
rect 106782 543910 106838 543966
rect 106906 543910 106962 543966
rect 107030 543910 107086 543966
rect 107154 543910 107210 543966
rect 68074 532272 68130 532328
rect 68198 532272 68254 532328
rect 68322 532272 68378 532328
rect 68446 532272 68502 532328
rect 68570 532272 68626 532328
rect 68694 532272 68750 532328
rect 68818 532272 68874 532328
rect 68942 532272 68998 532328
rect 69066 532272 69122 532328
rect 69190 532272 69246 532328
rect 69314 532272 69370 532328
rect 69438 532272 69494 532328
rect 69562 532272 69618 532328
rect 69686 532272 69742 532328
rect 69810 532272 69866 532328
rect 69934 532272 69990 532328
rect 70058 532272 70114 532328
rect 70182 532272 70238 532328
rect 70306 532272 70362 532328
rect 70430 532272 70486 532328
rect 70554 532272 70610 532328
rect 70678 532272 70734 532328
rect 70802 532272 70858 532328
rect 70926 532272 70982 532328
rect 71050 532272 71106 532328
rect 71174 532272 71230 532328
rect 71298 532272 71354 532328
rect 71422 532272 71478 532328
rect 71546 532272 71602 532328
rect 71670 532272 71726 532328
rect 71794 532272 71850 532328
rect 71918 532272 71974 532328
rect 72042 532272 72098 532328
rect 72166 532272 72222 532328
rect 72290 532272 72346 532328
rect 72414 532272 72470 532328
rect 72538 532272 72594 532328
rect 72662 532272 72718 532328
rect 72786 532272 72842 532328
rect 72910 532272 72966 532328
rect 73034 532272 73090 532328
rect 73158 532272 73214 532328
rect 73282 532272 73338 532328
rect 73406 532272 73462 532328
rect 73530 532272 73586 532328
rect 73654 532272 73710 532328
rect 73778 532272 73834 532328
rect 73902 532272 73958 532328
rect 74026 532272 74082 532328
rect 74150 532272 74206 532328
rect 74274 532272 74330 532328
rect 74398 532272 74454 532328
rect 74522 532272 74578 532328
rect 74646 532272 74702 532328
rect 74770 532272 74826 532328
rect 74894 532272 74950 532328
rect 75018 532272 75074 532328
rect 75142 532272 75198 532328
rect 75266 532272 75322 532328
rect 75390 532272 75446 532328
rect 84890 526272 84946 526328
rect 85014 526272 85070 526328
rect 85138 526272 85194 526328
rect 85262 526272 85318 526328
rect 85386 526272 85442 526328
rect 85510 526272 85566 526328
rect 85634 526272 85690 526328
rect 85758 526272 85814 526328
rect 85882 526272 85938 526328
rect 86006 526272 86062 526328
rect 86130 526272 86186 526328
rect 86254 526272 86310 526328
rect 86378 526272 86434 526328
rect 86502 526272 86558 526328
rect 86626 526272 86682 526328
rect 86750 526272 86806 526328
rect 86874 526272 86930 526328
rect 86998 526272 87054 526328
rect 87122 526272 87178 526328
rect 87246 526272 87302 526328
rect 87370 526272 87426 526328
rect 87494 526272 87550 526328
rect 87618 526272 87674 526328
rect 87742 526272 87798 526328
rect 87866 526272 87922 526328
rect 87990 526272 88046 526328
rect 88114 526272 88170 526328
rect 88238 526272 88294 526328
rect 88362 526272 88418 526328
rect 88486 526272 88542 526328
rect 88610 526272 88666 526328
rect 88734 526272 88790 526328
rect 88858 526272 88914 526328
rect 88982 526272 89038 526328
rect 89106 526272 89162 526328
rect 89230 526272 89286 526328
rect 89354 526272 89410 526328
rect 89478 526272 89534 526328
rect 89602 526272 89658 526328
rect 89726 526272 89782 526328
rect 89850 526272 89906 526328
rect 89974 526272 90030 526328
rect 90098 526272 90154 526328
rect 90222 526272 90278 526328
rect 90346 526272 90402 526328
rect 90470 526272 90526 526328
rect 90594 526272 90650 526328
rect 90718 526272 90774 526328
rect 90842 526272 90898 526328
rect 90966 526272 91022 526328
rect 91090 526272 91146 526328
rect 91214 526272 91270 526328
rect 91338 526272 91394 526328
rect 91462 526272 91518 526328
rect 91586 526272 91642 526328
rect 91710 526272 91766 526328
rect 91834 526272 91890 526328
rect 91958 526272 92014 526328
rect 92082 526272 92138 526328
rect 92206 526272 92262 526328
rect 92330 526272 92386 526328
rect 92454 526272 92510 526328
rect 92578 526272 92634 526328
rect 92702 526272 92758 526328
rect 92826 526272 92882 526328
rect 92950 526272 93006 526328
rect 93074 526272 93130 526328
rect 93198 526272 93254 526328
rect 93322 526272 93378 526328
rect 93446 526272 93502 526328
rect 93570 526272 93626 526328
rect 93694 526272 93750 526328
rect 93818 526272 93874 526328
rect 93942 526272 93998 526328
rect 94066 526272 94122 526328
rect 94190 526272 94246 526328
rect 94314 526272 94370 526328
rect 94438 526272 94494 526328
rect 94562 526272 94618 526328
rect 94686 526272 94742 526328
rect 94810 526272 94866 526328
rect 94934 526272 94990 526328
rect 95058 526272 95114 526328
rect 95182 526272 95238 526328
rect 95306 526272 95362 526328
rect 95430 526272 95486 526328
rect 95554 526272 95610 526328
rect 95678 526272 95734 526328
rect 95802 526272 95858 526328
rect 95926 526272 95982 526328
rect 96050 526272 96106 526328
rect 96174 526272 96230 526328
rect 96298 526272 96354 526328
rect 96422 526272 96478 526328
rect 96546 526272 96602 526328
rect 96670 526272 96726 526328
rect 96794 526272 96850 526328
rect 96918 526272 96974 526328
rect 97042 526272 97098 526328
rect 97166 526272 97222 526328
rect 97290 526272 97346 526328
rect 97414 526272 97470 526328
rect 97538 526272 97594 526328
rect 97662 526272 97718 526328
rect 97786 526272 97842 526328
rect 97910 526272 97966 526328
rect 98034 526272 98090 526328
rect 98158 526272 98214 526328
rect 98282 526272 98338 526328
rect 98406 526272 98462 526328
rect 98530 526272 98586 526328
rect 98654 526272 98710 526328
rect 84772 526034 84828 526090
rect 84896 526034 84952 526090
rect 85020 526034 85076 526090
rect 85144 526034 85200 526090
rect 85268 526034 85324 526090
rect 85392 526034 85448 526090
rect 85516 526034 85572 526090
rect 85640 526034 85696 526090
rect 85764 526034 85820 526090
rect 85888 526034 85944 526090
rect 86012 526034 86068 526090
rect 86136 526034 86192 526090
rect 86260 526034 86316 526090
rect 86384 526034 86440 526090
rect 86508 526034 86564 526090
rect 86632 526034 86688 526090
rect 86756 526034 86812 526090
rect 86880 526034 86936 526090
rect 87004 526034 87060 526090
rect 87128 526034 87184 526090
rect 87252 526034 87308 526090
rect 87376 526034 87432 526090
rect 87500 526034 87556 526090
rect 87624 526034 87680 526090
rect 87748 526034 87804 526090
rect 87872 526034 87928 526090
rect 87996 526034 88052 526090
rect 88120 526034 88176 526090
rect 88244 526034 88300 526090
rect 88368 526034 88424 526090
rect 88492 526034 88548 526090
rect 88616 526034 88672 526090
rect 88740 526034 88796 526090
rect 88864 526034 88920 526090
rect 88988 526034 89044 526090
rect 89112 526034 89168 526090
rect 89236 526034 89292 526090
rect 89360 526034 89416 526090
rect 89484 526034 89540 526090
rect 89608 526034 89664 526090
rect 89732 526034 89788 526090
rect 89856 526034 89912 526090
rect 89980 526034 90036 526090
rect 90104 526034 90160 526090
rect 90228 526034 90284 526090
rect 90352 526034 90408 526090
rect 90476 526034 90532 526090
rect 90600 526034 90656 526090
rect 90724 526034 90780 526090
rect 90848 526034 90904 526090
rect 90972 526034 91028 526090
rect 91096 526034 91152 526090
rect 91220 526034 91276 526090
rect 91344 526034 91400 526090
rect 91468 526034 91524 526090
rect 91592 526034 91648 526090
rect 91716 526034 91772 526090
rect 91840 526034 91896 526090
rect 91964 526034 92020 526090
rect 92088 526034 92144 526090
rect 92212 526034 92268 526090
rect 92336 526034 92392 526090
rect 92460 526034 92516 526090
rect 92584 526034 92640 526090
rect 92708 526034 92764 526090
rect 92832 526034 92888 526090
rect 92956 526034 93012 526090
rect 93080 526034 93136 526090
rect 93204 526034 93260 526090
rect 93328 526034 93384 526090
rect 93452 526034 93508 526090
rect 93576 526034 93632 526090
rect 93700 526034 93756 526090
rect 93824 526034 93880 526090
rect 93948 526034 94004 526090
rect 94072 526034 94128 526090
rect 94196 526034 94252 526090
rect 94320 526034 94376 526090
rect 94444 526034 94500 526090
rect 94568 526034 94624 526090
rect 94692 526034 94748 526090
rect 94816 526034 94872 526090
rect 94940 526034 94996 526090
rect 95064 526034 95120 526090
rect 95188 526034 95244 526090
rect 95312 526034 95368 526090
rect 95436 526034 95492 526090
rect 95560 526034 95616 526090
rect 95684 526034 95740 526090
rect 95808 526034 95864 526090
rect 95932 526034 95988 526090
rect 96056 526034 96112 526090
rect 96180 526034 96236 526090
rect 96304 526034 96360 526090
rect 96428 526034 96484 526090
rect 96552 526034 96608 526090
rect 96676 526034 96732 526090
rect 96800 526034 96856 526090
rect 96924 526034 96980 526090
rect 97048 526034 97104 526090
rect 97172 526034 97228 526090
rect 97296 526034 97352 526090
rect 97420 526034 97476 526090
rect 97544 526034 97600 526090
rect 97668 526034 97724 526090
rect 97792 526034 97848 526090
rect 97916 526034 97972 526090
rect 98040 526034 98096 526090
rect 98164 526034 98220 526090
rect 98288 526034 98344 526090
rect 98412 526034 98468 526090
rect 84772 525910 84828 525966
rect 84896 525910 84952 525966
rect 85020 525910 85076 525966
rect 85144 525910 85200 525966
rect 85268 525910 85324 525966
rect 85392 525910 85448 525966
rect 85516 525910 85572 525966
rect 85640 525910 85696 525966
rect 85764 525910 85820 525966
rect 85888 525910 85944 525966
rect 86012 525910 86068 525966
rect 86136 525910 86192 525966
rect 86260 525910 86316 525966
rect 86384 525910 86440 525966
rect 86508 525910 86564 525966
rect 86632 525910 86688 525966
rect 86756 525910 86812 525966
rect 86880 525910 86936 525966
rect 87004 525910 87060 525966
rect 87128 525910 87184 525966
rect 87252 525910 87308 525966
rect 87376 525910 87432 525966
rect 87500 525910 87556 525966
rect 87624 525910 87680 525966
rect 87748 525910 87804 525966
rect 87872 525910 87928 525966
rect 87996 525910 88052 525966
rect 88120 525910 88176 525966
rect 88244 525910 88300 525966
rect 88368 525910 88424 525966
rect 88492 525910 88548 525966
rect 88616 525910 88672 525966
rect 88740 525910 88796 525966
rect 88864 525910 88920 525966
rect 88988 525910 89044 525966
rect 89112 525910 89168 525966
rect 89236 525910 89292 525966
rect 89360 525910 89416 525966
rect 89484 525910 89540 525966
rect 89608 525910 89664 525966
rect 89732 525910 89788 525966
rect 89856 525910 89912 525966
rect 89980 525910 90036 525966
rect 90104 525910 90160 525966
rect 90228 525910 90284 525966
rect 90352 525910 90408 525966
rect 90476 525910 90532 525966
rect 90600 525910 90656 525966
rect 90724 525910 90780 525966
rect 90848 525910 90904 525966
rect 90972 525910 91028 525966
rect 91096 525910 91152 525966
rect 91220 525910 91276 525966
rect 91344 525910 91400 525966
rect 91468 525910 91524 525966
rect 91592 525910 91648 525966
rect 91716 525910 91772 525966
rect 91840 525910 91896 525966
rect 91964 525910 92020 525966
rect 92088 525910 92144 525966
rect 92212 525910 92268 525966
rect 92336 525910 92392 525966
rect 92460 525910 92516 525966
rect 92584 525910 92640 525966
rect 92708 525910 92764 525966
rect 92832 525910 92888 525966
rect 92956 525910 93012 525966
rect 93080 525910 93136 525966
rect 93204 525910 93260 525966
rect 93328 525910 93384 525966
rect 93452 525910 93508 525966
rect 93576 525910 93632 525966
rect 93700 525910 93756 525966
rect 93824 525910 93880 525966
rect 93948 525910 94004 525966
rect 94072 525910 94128 525966
rect 94196 525910 94252 525966
rect 94320 525910 94376 525966
rect 94444 525910 94500 525966
rect 94568 525910 94624 525966
rect 94692 525910 94748 525966
rect 94816 525910 94872 525966
rect 94940 525910 94996 525966
rect 95064 525910 95120 525966
rect 95188 525910 95244 525966
rect 95312 525910 95368 525966
rect 95436 525910 95492 525966
rect 95560 525910 95616 525966
rect 95684 525910 95740 525966
rect 95808 525910 95864 525966
rect 95932 525910 95988 525966
rect 96056 525910 96112 525966
rect 96180 525910 96236 525966
rect 96304 525910 96360 525966
rect 96428 525910 96484 525966
rect 96552 525910 96608 525966
rect 96676 525910 96732 525966
rect 96800 525910 96856 525966
rect 96924 525910 96980 525966
rect 97048 525910 97104 525966
rect 97172 525910 97228 525966
rect 97296 525910 97352 525966
rect 97420 525910 97476 525966
rect 97544 525910 97600 525966
rect 97668 525910 97724 525966
rect 97792 525910 97848 525966
rect 97916 525910 97972 525966
rect 98040 525910 98096 525966
rect 98164 525910 98220 525966
rect 98288 525910 98344 525966
rect 98412 525910 98468 525966
rect 60026 514356 60082 514412
rect 60150 514356 60206 514412
rect 60026 514232 60082 514288
rect 60150 514232 60206 514288
rect 60026 514108 60082 514164
rect 60150 514108 60206 514164
rect 60026 513984 60082 514040
rect 60150 513984 60206 514040
rect 60026 513860 60082 513916
rect 60150 513860 60206 513916
rect 60274 514356 60330 514412
rect 60398 514356 60454 514412
rect 60522 514356 60578 514412
rect 60646 514356 60702 514412
rect 60274 514232 60330 514288
rect 60398 514232 60454 514288
rect 60522 514232 60578 514288
rect 60646 514232 60702 514288
rect 60274 514108 60330 514164
rect 60398 514108 60454 514164
rect 60522 514108 60578 514164
rect 60646 514108 60702 514164
rect 60274 513984 60330 514040
rect 60398 513984 60454 514040
rect 60522 513984 60578 514040
rect 60646 513984 60702 514040
rect 60274 513860 60330 513916
rect 60398 513860 60454 513916
rect 60522 513860 60578 513916
rect 60646 513860 60702 513916
rect 60770 514356 60826 514412
rect 60894 514356 60950 514412
rect 61018 514356 61074 514412
rect 61142 514356 61198 514412
rect 60770 514232 60826 514288
rect 60894 514232 60950 514288
rect 61018 514232 61074 514288
rect 61142 514232 61198 514288
rect 60770 514108 60826 514164
rect 60894 514108 60950 514164
rect 61018 514108 61074 514164
rect 61142 514108 61198 514164
rect 60770 513984 60826 514040
rect 60894 513984 60950 514040
rect 61018 513984 61074 514040
rect 61142 513984 61198 514040
rect 60770 513860 60826 513916
rect 60894 513860 60950 513916
rect 61018 513860 61074 513916
rect 61142 513860 61198 513916
rect 61266 514356 61322 514412
rect 61390 514356 61446 514412
rect 61514 514356 61570 514412
rect 61638 514356 61694 514412
rect 61266 514232 61322 514288
rect 61390 514232 61446 514288
rect 61514 514232 61570 514288
rect 61638 514232 61694 514288
rect 61266 514108 61322 514164
rect 61390 514108 61446 514164
rect 61514 514108 61570 514164
rect 61638 514108 61694 514164
rect 61266 513984 61322 514040
rect 61390 513984 61446 514040
rect 61514 513984 61570 514040
rect 61638 513984 61694 514040
rect 61266 513860 61322 513916
rect 61390 513860 61446 513916
rect 61514 513860 61570 513916
rect 61638 513860 61694 513916
rect 61762 514356 61818 514412
rect 61886 514356 61942 514412
rect 62010 514356 62066 514412
rect 62134 514356 62190 514412
rect 61762 514232 61818 514288
rect 61886 514232 61942 514288
rect 62010 514232 62066 514288
rect 62134 514232 62190 514288
rect 61762 514108 61818 514164
rect 61886 514108 61942 514164
rect 62010 514108 62066 514164
rect 62134 514108 62190 514164
rect 61762 513984 61818 514040
rect 61886 513984 61942 514040
rect 62010 513984 62066 514040
rect 62134 513984 62190 514040
rect 61762 513860 61818 513916
rect 61886 513860 61942 513916
rect 62010 513860 62066 513916
rect 62134 513860 62190 513916
rect 62258 514356 62314 514412
rect 62382 514356 62438 514412
rect 62506 514356 62562 514412
rect 62630 514356 62686 514412
rect 62258 514232 62314 514288
rect 62382 514232 62438 514288
rect 62506 514232 62562 514288
rect 62630 514232 62686 514288
rect 62258 514108 62314 514164
rect 62382 514108 62438 514164
rect 62506 514108 62562 514164
rect 62630 514108 62686 514164
rect 62258 513984 62314 514040
rect 62382 513984 62438 514040
rect 62506 513984 62562 514040
rect 62630 513984 62686 514040
rect 62258 513860 62314 513916
rect 62382 513860 62438 513916
rect 62506 513860 62562 513916
rect 62630 513860 62686 513916
rect 62754 514356 62810 514412
rect 62878 514356 62934 514412
rect 63002 514356 63058 514412
rect 63126 514356 63182 514412
rect 62754 514232 62810 514288
rect 62878 514232 62934 514288
rect 63002 514232 63058 514288
rect 63126 514232 63182 514288
rect 62754 514108 62810 514164
rect 62878 514108 62934 514164
rect 63002 514108 63058 514164
rect 63126 514108 63182 514164
rect 62754 513984 62810 514040
rect 62878 513984 62934 514040
rect 63002 513984 63058 514040
rect 63126 513984 63182 514040
rect 62754 513860 62810 513916
rect 62878 513860 62934 513916
rect 63002 513860 63058 513916
rect 63126 513860 63182 513916
rect 63250 514356 63306 514412
rect 63374 514356 63430 514412
rect 63498 514356 63554 514412
rect 63622 514356 63678 514412
rect 63250 514232 63306 514288
rect 63374 514232 63430 514288
rect 63498 514232 63554 514288
rect 63622 514232 63678 514288
rect 63250 514108 63306 514164
rect 63374 514108 63430 514164
rect 63498 514108 63554 514164
rect 63622 514108 63678 514164
rect 63250 513984 63306 514040
rect 63374 513984 63430 514040
rect 63498 513984 63554 514040
rect 63622 513984 63678 514040
rect 63250 513860 63306 513916
rect 63374 513860 63430 513916
rect 63498 513860 63554 513916
rect 63622 513860 63678 513916
rect 63746 514356 63802 514412
rect 63870 514356 63926 514412
rect 63994 514356 64050 514412
rect 64118 514356 64174 514412
rect 63746 514232 63802 514288
rect 63870 514232 63926 514288
rect 63994 514232 64050 514288
rect 64118 514232 64174 514288
rect 63746 514108 63802 514164
rect 63870 514108 63926 514164
rect 63994 514108 64050 514164
rect 64118 514108 64174 514164
rect 63746 513984 63802 514040
rect 63870 513984 63926 514040
rect 63994 513984 64050 514040
rect 64118 513984 64174 514040
rect 63746 513860 63802 513916
rect 63870 513860 63926 513916
rect 63994 513860 64050 513916
rect 64118 513860 64174 513916
rect 78970 508375 79026 508431
rect 79094 508375 79150 508431
rect 79218 508375 79274 508431
rect 79342 508375 79398 508431
rect 79466 508375 79522 508431
rect 79590 508375 79646 508431
rect 79714 508375 79770 508431
rect 79838 508375 79894 508431
rect 79962 508375 80018 508431
rect 80086 508375 80142 508431
rect 80210 508375 80266 508431
rect 80334 508375 80390 508431
rect 80458 508375 80514 508431
rect 80582 508375 80638 508431
rect 80706 508375 80762 508431
rect 80830 508375 80886 508431
rect 80954 508375 81010 508431
rect 81078 508375 81134 508431
rect 81202 508375 81258 508431
rect 81326 508375 81382 508431
rect 81450 508375 81506 508431
rect 81574 508375 81630 508431
rect 81698 508375 81754 508431
rect 81822 508375 81878 508431
rect 81946 508375 82002 508431
rect 82070 508375 82126 508431
rect 82194 508375 82250 508431
rect 82318 508375 82374 508431
rect 82442 508375 82498 508431
rect 82566 508375 82622 508431
rect 82690 508375 82746 508431
rect 82814 508375 82870 508431
rect 82938 508375 82994 508431
rect 83062 508375 83118 508431
rect 83186 508375 83242 508431
rect 83310 508375 83366 508431
rect 83434 508375 83490 508431
rect 83558 508375 83614 508431
rect 83682 508375 83738 508431
rect 83806 508375 83862 508431
rect 83930 508375 83986 508431
rect 84054 508375 84110 508431
rect 78850 508152 78906 508208
rect 78974 508152 79030 508208
rect 79098 508152 79154 508208
rect 79222 508152 79278 508208
rect 79346 508152 79402 508208
rect 79470 508152 79526 508208
rect 79594 508152 79650 508208
rect 79718 508152 79774 508208
rect 79842 508152 79898 508208
rect 79966 508152 80022 508208
rect 80090 508152 80146 508208
rect 80214 508152 80270 508208
rect 80338 508152 80394 508208
rect 80462 508152 80518 508208
rect 80586 508152 80642 508208
rect 80710 508152 80766 508208
rect 80834 508152 80890 508208
rect 80958 508152 81014 508208
rect 81082 508152 81138 508208
rect 81206 508152 81262 508208
rect 81330 508152 81386 508208
rect 81454 508152 81510 508208
rect 81578 508152 81634 508208
rect 81702 508152 81758 508208
rect 81826 508152 81882 508208
rect 81950 508152 82006 508208
rect 82074 508152 82130 508208
rect 82198 508152 82254 508208
rect 82322 508152 82378 508208
rect 82446 508152 82502 508208
rect 82570 508152 82626 508208
rect 82694 508152 82750 508208
rect 82818 508152 82874 508208
rect 82942 508152 82998 508208
rect 83066 508152 83122 508208
rect 83190 508152 83246 508208
rect 83314 508152 83370 508208
rect 83438 508152 83494 508208
rect 83562 508152 83618 508208
rect 83686 508152 83742 508208
rect 83810 508152 83866 508208
rect 83934 508152 83990 508208
rect 67964 496272 68020 496328
rect 68088 496272 68144 496328
rect 68212 496272 68268 496328
rect 68336 496272 68392 496328
rect 68460 496272 68516 496328
rect 68584 496272 68640 496328
rect 68708 496272 68764 496328
rect 68832 496272 68888 496328
rect 68956 496272 69012 496328
rect 69080 496272 69136 496328
rect 69204 496272 69260 496328
rect 69328 496272 69384 496328
rect 69452 496272 69508 496328
rect 69576 496272 69632 496328
rect 69700 496272 69756 496328
rect 69824 496272 69880 496328
rect 69948 496272 70004 496328
rect 70072 496272 70128 496328
rect 70196 496272 70252 496328
rect 70320 496272 70376 496328
rect 70444 496272 70500 496328
rect 70568 496272 70624 496328
rect 70692 496272 70748 496328
rect 70816 496272 70872 496328
rect 70940 496272 70996 496328
rect 71064 496272 71120 496328
rect 71188 496272 71244 496328
rect 71312 496272 71368 496328
rect 71436 496272 71492 496328
rect 71560 496272 71616 496328
rect 71684 496272 71740 496328
rect 71808 496272 71864 496328
rect 71932 496272 71988 496328
rect 72056 496272 72112 496328
rect 72180 496272 72236 496328
rect 72304 496272 72360 496328
rect 72428 496272 72484 496328
rect 72552 496272 72608 496328
rect 72676 496272 72732 496328
rect 72800 496272 72856 496328
rect 72924 496272 72980 496328
rect 73048 496272 73104 496328
rect 73172 496272 73228 496328
rect 73296 496272 73352 496328
rect 73420 496272 73476 496328
rect 73544 496272 73600 496328
rect 73668 496272 73724 496328
rect 73792 496272 73848 496328
rect 73916 496272 73972 496328
rect 74040 496272 74096 496328
rect 74164 496272 74220 496328
rect 74288 496272 74344 496328
rect 74412 496272 74468 496328
rect 74536 496272 74592 496328
rect 74660 496272 74716 496328
rect 68208 496032 68264 496088
rect 68332 496032 68388 496088
rect 68456 496032 68512 496088
rect 68580 496032 68636 496088
rect 68704 496032 68760 496088
rect 68828 496032 68884 496088
rect 68952 496032 69008 496088
rect 69076 496032 69132 496088
rect 69200 496032 69256 496088
rect 69324 496032 69380 496088
rect 69448 496032 69504 496088
rect 69572 496032 69628 496088
rect 69696 496032 69752 496088
rect 69820 496032 69876 496088
rect 69944 496032 70000 496088
rect 70068 496032 70124 496088
rect 70192 496032 70248 496088
rect 70316 496032 70372 496088
rect 70440 496032 70496 496088
rect 70564 496032 70620 496088
rect 70688 496032 70744 496088
rect 70812 496032 70868 496088
rect 70936 496032 70992 496088
rect 71060 496032 71116 496088
rect 71184 496032 71240 496088
rect 71308 496032 71364 496088
rect 71432 496032 71488 496088
rect 71556 496032 71612 496088
rect 71680 496032 71736 496088
rect 71804 496032 71860 496088
rect 71928 496032 71984 496088
rect 72052 496032 72108 496088
rect 72176 496032 72232 496088
rect 72300 496032 72356 496088
rect 72424 496032 72480 496088
rect 72548 496032 72604 496088
rect 72672 496032 72728 496088
rect 72796 496032 72852 496088
rect 72920 496032 72976 496088
rect 73044 496032 73100 496088
rect 73168 496032 73224 496088
rect 73292 496032 73348 496088
rect 73416 496032 73472 496088
rect 73540 496032 73596 496088
rect 73664 496032 73720 496088
rect 73788 496032 73844 496088
rect 73912 496032 73968 496088
rect 74036 496032 74092 496088
rect 74160 496032 74216 496088
rect 74284 496032 74340 496088
rect 74408 496032 74464 496088
rect 74532 496032 74588 496088
rect 74656 496032 74712 496088
rect 66954 490294 67010 490350
rect 67078 490294 67134 490350
rect 67202 490294 67258 490350
rect 67326 490294 67382 490350
rect 66954 490170 67010 490226
rect 67078 490170 67134 490226
rect 67202 490170 67258 490226
rect 67326 490170 67382 490226
rect 66954 490046 67010 490102
rect 67078 490046 67134 490102
rect 67202 490046 67258 490102
rect 67326 490046 67382 490102
rect 66954 489922 67010 489978
rect 67078 489922 67134 489978
rect 67202 489922 67258 489978
rect 67326 489922 67382 489978
rect 60172 409742 60228 409798
rect 60284 408122 60340 408178
rect 60508 404740 60564 404758
rect 60508 404702 60564 404740
rect 60284 383102 60340 383158
rect 60172 374642 60228 374698
rect 57932 301742 57988 301798
rect 56924 297062 56980 297118
rect 58156 295622 58212 295678
rect 60172 368162 60228 368218
rect 58492 296702 58548 296758
rect 58716 295442 58772 295498
rect 60508 350028 60564 350038
rect 60508 349982 60564 350028
rect 60172 335942 60228 335998
rect 60172 329282 60228 329338
rect 60508 344428 60564 344458
rect 60508 344402 60564 344428
rect 60396 324268 60452 324298
rect 60396 324242 60452 324268
rect 60508 301562 60564 301618
rect 60284 288782 60340 288838
rect 60172 286982 60228 287038
rect 60060 283562 60116 283618
rect 58604 281942 58660 281998
rect 60732 374822 60788 374878
rect 60732 368004 60788 368038
rect 60732 367982 60788 368004
rect 60732 366362 60788 366418
rect 60732 335762 60788 335818
rect 60732 326762 60788 326818
rect 60732 307524 60788 307558
rect 60732 307502 60788 307524
rect 66954 472294 67010 472350
rect 67078 472294 67134 472350
rect 67202 472294 67258 472350
rect 67326 472294 67382 472350
rect 66954 472170 67010 472226
rect 67078 472170 67134 472226
rect 67202 472170 67258 472226
rect 67326 472170 67382 472226
rect 66954 472046 67010 472102
rect 67078 472046 67134 472102
rect 67202 472046 67258 472102
rect 67326 472046 67382 472102
rect 66954 471922 67010 471978
rect 67078 471922 67134 471978
rect 67202 471922 67258 471978
rect 67326 471922 67382 471978
rect 66954 454294 67010 454350
rect 67078 454294 67134 454350
rect 67202 454294 67258 454350
rect 67326 454294 67382 454350
rect 66954 454170 67010 454226
rect 67078 454170 67134 454226
rect 67202 454170 67258 454226
rect 67326 454170 67382 454226
rect 66954 454046 67010 454102
rect 67078 454046 67134 454102
rect 67202 454046 67258 454102
rect 67326 454046 67382 454102
rect 66954 453922 67010 453978
rect 67078 453922 67134 453978
rect 67202 453922 67258 453978
rect 67326 453922 67382 453978
rect 66954 436294 67010 436350
rect 67078 436294 67134 436350
rect 67202 436294 67258 436350
rect 67326 436294 67382 436350
rect 66954 436170 67010 436226
rect 67078 436170 67134 436226
rect 67202 436170 67258 436226
rect 67326 436170 67382 436226
rect 66954 436046 67010 436102
rect 67078 436046 67134 436102
rect 67202 436046 67258 436102
rect 67326 436046 67382 436102
rect 66954 435922 67010 435978
rect 67078 435922 67134 435978
rect 67202 435922 67258 435978
rect 67326 435922 67382 435978
rect 64518 418294 64574 418350
rect 64642 418294 64698 418350
rect 64518 418170 64574 418226
rect 64642 418170 64698 418226
rect 64518 418046 64574 418102
rect 64642 418046 64698 418102
rect 64518 417922 64574 417978
rect 64642 417922 64698 417978
rect 64518 400294 64574 400350
rect 64642 400294 64698 400350
rect 64518 400170 64574 400226
rect 64642 400170 64698 400226
rect 64518 400046 64574 400102
rect 64642 400046 64698 400102
rect 64518 399922 64574 399978
rect 64642 399922 64698 399978
rect 64518 382294 64574 382350
rect 64642 382294 64698 382350
rect 64518 382170 64574 382226
rect 64642 382170 64698 382226
rect 64518 382046 64574 382102
rect 64642 382046 64698 382102
rect 64518 381922 64574 381978
rect 64642 381922 64698 381978
rect 64518 364294 64574 364350
rect 64642 364294 64698 364350
rect 64518 364170 64574 364226
rect 64642 364170 64698 364226
rect 64518 364046 64574 364102
rect 64642 364046 64698 364102
rect 64518 363922 64574 363978
rect 64642 363922 64698 363978
rect 64518 346294 64574 346350
rect 64642 346294 64698 346350
rect 64518 346170 64574 346226
rect 64642 346170 64698 346226
rect 64518 346046 64574 346102
rect 64642 346046 64698 346102
rect 64518 345922 64574 345978
rect 64642 345922 64698 345978
rect 64518 328294 64574 328350
rect 64642 328294 64698 328350
rect 64518 328170 64574 328226
rect 64642 328170 64698 328226
rect 64518 328046 64574 328102
rect 64642 328046 64698 328102
rect 64518 327922 64574 327978
rect 64642 327922 64698 327978
rect 64518 310294 64574 310350
rect 64642 310294 64698 310350
rect 64518 310170 64574 310226
rect 64642 310170 64698 310226
rect 64518 310046 64574 310102
rect 64642 310046 64698 310102
rect 64518 309922 64574 309978
rect 64642 309922 64698 309978
rect 70674 478294 70730 478350
rect 70798 478294 70854 478350
rect 70922 478294 70978 478350
rect 71046 478294 71102 478350
rect 70674 478170 70730 478226
rect 70798 478170 70854 478226
rect 70922 478170 70978 478226
rect 71046 478170 71102 478226
rect 70674 478046 70730 478102
rect 70798 478046 70854 478102
rect 70922 478046 70978 478102
rect 71046 478046 71102 478102
rect 70674 477922 70730 477978
rect 70798 477922 70854 477978
rect 70922 477922 70978 477978
rect 71046 477922 71102 477978
rect 70674 460294 70730 460350
rect 70798 460294 70854 460350
rect 70922 460294 70978 460350
rect 71046 460294 71102 460350
rect 70674 460170 70730 460226
rect 70798 460170 70854 460226
rect 70922 460170 70978 460226
rect 71046 460170 71102 460226
rect 70674 460046 70730 460102
rect 70798 460046 70854 460102
rect 70922 460046 70978 460102
rect 71046 460046 71102 460102
rect 70674 459922 70730 459978
rect 70798 459922 70854 459978
rect 70922 459922 70978 459978
rect 71046 459922 71102 459978
rect 70674 442294 70730 442350
rect 70798 442294 70854 442350
rect 70922 442294 70978 442350
rect 71046 442294 71102 442350
rect 70674 442170 70730 442226
rect 70798 442170 70854 442226
rect 70922 442170 70978 442226
rect 71046 442170 71102 442226
rect 70674 442046 70730 442102
rect 70798 442046 70854 442102
rect 70922 442046 70978 442102
rect 71046 442046 71102 442102
rect 70674 441922 70730 441978
rect 70798 441922 70854 441978
rect 70922 441922 70978 441978
rect 71046 441922 71102 441978
rect 69468 430982 69524 431038
rect 66954 418294 67010 418350
rect 67078 418294 67134 418350
rect 67202 418294 67258 418350
rect 67326 418294 67382 418350
rect 66954 418170 67010 418226
rect 67078 418170 67134 418226
rect 67202 418170 67258 418226
rect 67326 418170 67382 418226
rect 66954 418046 67010 418102
rect 67078 418046 67134 418102
rect 67202 418046 67258 418102
rect 67326 418046 67382 418102
rect 66954 417922 67010 417978
rect 67078 417922 67134 417978
rect 67202 417922 67258 417978
rect 67326 417922 67382 417978
rect 66954 400294 67010 400350
rect 67078 400294 67134 400350
rect 67202 400294 67258 400350
rect 67326 400294 67382 400350
rect 66954 400170 67010 400226
rect 67078 400170 67134 400226
rect 67202 400170 67258 400226
rect 67326 400170 67382 400226
rect 66954 400046 67010 400102
rect 67078 400046 67134 400102
rect 67202 400046 67258 400102
rect 67326 400046 67382 400102
rect 66954 399922 67010 399978
rect 67078 399922 67134 399978
rect 67202 399922 67258 399978
rect 67326 399922 67382 399978
rect 66954 382294 67010 382350
rect 67078 382294 67134 382350
rect 67202 382294 67258 382350
rect 67326 382294 67382 382350
rect 66954 382170 67010 382226
rect 67078 382170 67134 382226
rect 67202 382170 67258 382226
rect 67326 382170 67382 382226
rect 66954 382046 67010 382102
rect 67078 382046 67134 382102
rect 67202 382046 67258 382102
rect 67326 382046 67382 382102
rect 66954 381922 67010 381978
rect 67078 381922 67134 381978
rect 67202 381922 67258 381978
rect 67326 381922 67382 381978
rect 66954 364294 67010 364350
rect 67078 364294 67134 364350
rect 67202 364294 67258 364350
rect 67326 364294 67382 364350
rect 66954 364170 67010 364226
rect 67078 364170 67134 364226
rect 67202 364170 67258 364226
rect 67326 364170 67382 364226
rect 66954 364046 67010 364102
rect 67078 364046 67134 364102
rect 67202 364046 67258 364102
rect 67326 364046 67382 364102
rect 66954 363922 67010 363978
rect 67078 363922 67134 363978
rect 67202 363922 67258 363978
rect 67326 363922 67382 363978
rect 97674 490294 97730 490350
rect 97798 490294 97854 490350
rect 97922 490294 97978 490350
rect 98046 490294 98102 490350
rect 97674 490170 97730 490226
rect 97798 490170 97854 490226
rect 97922 490170 97978 490226
rect 98046 490170 98102 490226
rect 97674 490046 97730 490102
rect 97798 490046 97854 490102
rect 97922 490046 97978 490102
rect 98046 490046 98102 490102
rect 97674 489922 97730 489978
rect 97798 489922 97854 489978
rect 97922 489922 97978 489978
rect 98046 489922 98102 489978
rect 97674 472294 97730 472350
rect 97798 472294 97854 472350
rect 97922 472294 97978 472350
rect 98046 472294 98102 472350
rect 97674 472170 97730 472226
rect 97798 472170 97854 472226
rect 97922 472170 97978 472226
rect 98046 472170 98102 472226
rect 97674 472046 97730 472102
rect 97798 472046 97854 472102
rect 97922 472046 97978 472102
rect 98046 472046 98102 472102
rect 97674 471922 97730 471978
rect 97798 471922 97854 471978
rect 97922 471922 97978 471978
rect 98046 471922 98102 471978
rect 97674 454294 97730 454350
rect 97798 454294 97854 454350
rect 97922 454294 97978 454350
rect 98046 454294 98102 454350
rect 97674 454170 97730 454226
rect 97798 454170 97854 454226
rect 97922 454170 97978 454226
rect 98046 454170 98102 454226
rect 97674 454046 97730 454102
rect 97798 454046 97854 454102
rect 97922 454046 97978 454102
rect 98046 454046 98102 454102
rect 97674 453922 97730 453978
rect 97798 453922 97854 453978
rect 97922 453922 97978 453978
rect 98046 453922 98102 453978
rect 97674 436294 97730 436350
rect 97798 436294 97854 436350
rect 97922 436294 97978 436350
rect 98046 436294 98102 436350
rect 97674 436170 97730 436226
rect 97798 436170 97854 436226
rect 97922 436170 97978 436226
rect 98046 436170 98102 436226
rect 97674 436046 97730 436102
rect 97798 436046 97854 436102
rect 97922 436046 97978 436102
rect 98046 436046 98102 436102
rect 97674 435922 97730 435978
rect 97798 435922 97854 435978
rect 97922 435922 97978 435978
rect 98046 435922 98102 435978
rect 74844 429380 74900 429418
rect 74844 429362 74900 429380
rect 70674 424294 70730 424350
rect 70798 424294 70854 424350
rect 70922 424294 70978 424350
rect 71046 424294 71102 424350
rect 70674 424170 70730 424226
rect 70798 424170 70854 424226
rect 70922 424170 70978 424226
rect 71046 424170 71102 424226
rect 70674 424046 70730 424102
rect 70798 424046 70854 424102
rect 70922 424046 70978 424102
rect 71046 424046 71102 424102
rect 70674 423922 70730 423978
rect 70798 423922 70854 423978
rect 70922 423922 70978 423978
rect 71046 423922 71102 423978
rect 70674 406294 70730 406350
rect 70798 406294 70854 406350
rect 70922 406294 70978 406350
rect 71046 406294 71102 406350
rect 70674 406170 70730 406226
rect 70798 406170 70854 406226
rect 70922 406170 70978 406226
rect 71046 406170 71102 406226
rect 70674 406046 70730 406102
rect 70798 406046 70854 406102
rect 70922 406046 70978 406102
rect 71046 406046 71102 406102
rect 70674 405922 70730 405978
rect 70798 405922 70854 405978
rect 70922 405922 70978 405978
rect 71046 405922 71102 405978
rect 70674 388294 70730 388350
rect 70798 388294 70854 388350
rect 70922 388294 70978 388350
rect 71046 388294 71102 388350
rect 70674 388170 70730 388226
rect 70798 388170 70854 388226
rect 70922 388170 70978 388226
rect 71046 388170 71102 388226
rect 70674 388046 70730 388102
rect 70798 388046 70854 388102
rect 70922 388046 70978 388102
rect 71046 388046 71102 388102
rect 70674 387922 70730 387978
rect 70798 387922 70854 387978
rect 70922 387922 70978 387978
rect 71046 387922 71102 387978
rect 70674 370294 70730 370350
rect 70798 370294 70854 370350
rect 70922 370294 70978 370350
rect 71046 370294 71102 370350
rect 70674 370170 70730 370226
rect 70798 370170 70854 370226
rect 70922 370170 70978 370226
rect 71046 370170 71102 370226
rect 70674 370046 70730 370102
rect 70798 370046 70854 370102
rect 70922 370046 70978 370102
rect 71046 370046 71102 370102
rect 70674 369922 70730 369978
rect 70798 369922 70854 369978
rect 70922 369922 70978 369978
rect 71046 369922 71102 369978
rect 70674 352294 70730 352350
rect 70798 352294 70854 352350
rect 70922 352294 70978 352350
rect 71046 352294 71102 352350
rect 70674 352170 70730 352226
rect 70798 352170 70854 352226
rect 70922 352170 70978 352226
rect 71046 352170 71102 352226
rect 70674 352046 70730 352102
rect 70798 352046 70854 352102
rect 70922 352046 70978 352102
rect 71046 352046 71102 352102
rect 70674 351922 70730 351978
rect 70798 351922 70854 351978
rect 70922 351922 70978 351978
rect 71046 351922 71102 351978
rect 66954 346294 67010 346350
rect 67078 346294 67134 346350
rect 67202 346294 67258 346350
rect 67326 346294 67382 346350
rect 66954 346170 67010 346226
rect 67078 346170 67134 346226
rect 67202 346170 67258 346226
rect 67326 346170 67382 346226
rect 66954 346046 67010 346102
rect 67078 346046 67134 346102
rect 67202 346046 67258 346102
rect 67326 346046 67382 346102
rect 66954 345922 67010 345978
rect 67078 345922 67134 345978
rect 67202 345922 67258 345978
rect 67326 345922 67382 345978
rect 66954 328294 67010 328350
rect 67078 328294 67134 328350
rect 67202 328294 67258 328350
rect 67326 328294 67382 328350
rect 66954 328170 67010 328226
rect 67078 328170 67134 328226
rect 67202 328170 67258 328226
rect 67326 328170 67382 328226
rect 66954 328046 67010 328102
rect 67078 328046 67134 328102
rect 67202 328046 67258 328102
rect 67326 328046 67382 328102
rect 66954 327922 67010 327978
rect 67078 327922 67134 327978
rect 67202 327922 67258 327978
rect 67326 327922 67382 327978
rect 66954 310294 67010 310350
rect 67078 310294 67134 310350
rect 67202 310294 67258 310350
rect 67326 310294 67382 310350
rect 66954 310170 67010 310226
rect 67078 310170 67134 310226
rect 67202 310170 67258 310226
rect 67326 310170 67382 310226
rect 66954 310046 67010 310102
rect 67078 310046 67134 310102
rect 67202 310046 67258 310102
rect 67326 310046 67382 310102
rect 66954 309922 67010 309978
rect 67078 309922 67134 309978
rect 67202 309922 67258 309978
rect 67326 309922 67382 309978
rect 66954 292294 67010 292350
rect 67078 292294 67134 292350
rect 67202 292294 67258 292350
rect 67326 292294 67382 292350
rect 66954 292170 67010 292226
rect 67078 292170 67134 292226
rect 67202 292170 67258 292226
rect 67326 292170 67382 292226
rect 66954 292046 67010 292102
rect 67078 292046 67134 292102
rect 67202 292046 67258 292102
rect 67326 292046 67382 292102
rect 66954 291922 67010 291978
rect 67078 291922 67134 291978
rect 67202 291922 67258 291978
rect 67326 291922 67382 291978
rect 69692 349982 69748 350038
rect 69692 290402 69748 290458
rect 70674 334294 70730 334350
rect 70798 334294 70854 334350
rect 70922 334294 70978 334350
rect 71046 334294 71102 334350
rect 70674 334170 70730 334226
rect 70798 334170 70854 334226
rect 70922 334170 70978 334226
rect 71046 334170 71102 334226
rect 70674 334046 70730 334102
rect 70798 334046 70854 334102
rect 70922 334046 70978 334102
rect 71046 334046 71102 334102
rect 70674 333922 70730 333978
rect 70798 333922 70854 333978
rect 70922 333922 70978 333978
rect 71046 333922 71102 333978
rect 74732 326762 74788 326818
rect 70674 316294 70730 316350
rect 70798 316294 70854 316350
rect 70922 316294 70978 316350
rect 71046 316294 71102 316350
rect 70674 316170 70730 316226
rect 70798 316170 70854 316226
rect 70922 316170 70978 316226
rect 71046 316170 71102 316226
rect 70674 316046 70730 316102
rect 70798 316046 70854 316102
rect 70922 316046 70978 316102
rect 71046 316046 71102 316102
rect 70674 315922 70730 315978
rect 70798 315922 70854 315978
rect 70922 315922 70978 315978
rect 71046 315922 71102 315978
rect 70674 298294 70730 298350
rect 70798 298294 70854 298350
rect 70922 298294 70978 298350
rect 71046 298294 71102 298350
rect 70674 298170 70730 298226
rect 70798 298170 70854 298226
rect 70922 298170 70978 298226
rect 71046 298170 71102 298226
rect 70674 298046 70730 298102
rect 70798 298046 70854 298102
rect 70922 298046 70978 298102
rect 71046 298046 71102 298102
rect 70674 297922 70730 297978
rect 70798 297922 70854 297978
rect 70922 297922 70978 297978
rect 71046 297922 71102 297978
rect 66954 274294 67010 274350
rect 67078 274294 67134 274350
rect 67202 274294 67258 274350
rect 67326 274294 67382 274350
rect 66954 274170 67010 274226
rect 67078 274170 67134 274226
rect 67202 274170 67258 274226
rect 67326 274170 67382 274226
rect 66954 274046 67010 274102
rect 67078 274046 67134 274102
rect 67202 274046 67258 274102
rect 67326 274046 67382 274102
rect 66954 273922 67010 273978
rect 67078 273922 67134 273978
rect 67202 273922 67258 273978
rect 67326 273922 67382 273978
rect 66954 256294 67010 256350
rect 67078 256294 67134 256350
rect 67202 256294 67258 256350
rect 67326 256294 67382 256350
rect 66954 256170 67010 256226
rect 67078 256170 67134 256226
rect 67202 256170 67258 256226
rect 67326 256170 67382 256226
rect 66954 256046 67010 256102
rect 67078 256046 67134 256102
rect 67202 256046 67258 256102
rect 67326 256046 67382 256102
rect 66954 255922 67010 255978
rect 67078 255922 67134 255978
rect 67202 255922 67258 255978
rect 67326 255922 67382 255978
rect 66954 238294 67010 238350
rect 67078 238294 67134 238350
rect 67202 238294 67258 238350
rect 67326 238294 67382 238350
rect 66954 238170 67010 238226
rect 67078 238170 67134 238226
rect 67202 238170 67258 238226
rect 67326 238170 67382 238226
rect 66954 238046 67010 238102
rect 67078 238046 67134 238102
rect 67202 238046 67258 238102
rect 67326 238046 67382 238102
rect 66954 237922 67010 237978
rect 67078 237922 67134 237978
rect 67202 237922 67258 237978
rect 67326 237922 67382 237978
rect 70674 280294 70730 280350
rect 70798 280294 70854 280350
rect 70922 280294 70978 280350
rect 71046 280294 71102 280350
rect 70674 280170 70730 280226
rect 70798 280170 70854 280226
rect 70922 280170 70978 280226
rect 71046 280170 71102 280226
rect 70674 280046 70730 280102
rect 70798 280046 70854 280102
rect 70922 280046 70978 280102
rect 71046 280046 71102 280102
rect 70674 279922 70730 279978
rect 70798 279922 70854 279978
rect 70922 279922 70978 279978
rect 71046 279922 71102 279978
rect 70674 262294 70730 262350
rect 70798 262294 70854 262350
rect 70922 262294 70978 262350
rect 71046 262294 71102 262350
rect 70674 262170 70730 262226
rect 70798 262170 70854 262226
rect 70922 262170 70978 262226
rect 71046 262170 71102 262226
rect 70674 262046 70730 262102
rect 70798 262046 70854 262102
rect 70922 262046 70978 262102
rect 71046 262046 71102 262102
rect 70674 261922 70730 261978
rect 70798 261922 70854 261978
rect 70922 261922 70978 261978
rect 71046 261922 71102 261978
rect 73052 324242 73108 324298
rect 82908 432062 82964 432118
rect 77532 431882 77588 431938
rect 80220 428462 80276 428518
rect 79878 424294 79934 424350
rect 80002 424294 80058 424350
rect 79878 424170 79934 424226
rect 80002 424170 80058 424226
rect 79878 424046 79934 424102
rect 80002 424046 80058 424102
rect 79878 423922 79934 423978
rect 80002 423922 80058 423978
rect 79878 406294 79934 406350
rect 80002 406294 80058 406350
rect 79878 406170 79934 406226
rect 80002 406170 80058 406226
rect 79878 406046 79934 406102
rect 80002 406046 80058 406102
rect 79878 405922 79934 405978
rect 80002 405922 80058 405978
rect 79878 388294 79934 388350
rect 80002 388294 80058 388350
rect 79878 388170 79934 388226
rect 80002 388170 80058 388226
rect 79878 388046 79934 388102
rect 80002 388046 80058 388102
rect 79878 387922 79934 387978
rect 80002 387922 80058 387978
rect 79878 370294 79934 370350
rect 80002 370294 80058 370350
rect 79878 370170 79934 370226
rect 80002 370170 80058 370226
rect 79878 370046 79934 370102
rect 80002 370046 80058 370102
rect 79878 369922 79934 369978
rect 80002 369922 80058 369978
rect 79878 352294 79934 352350
rect 80002 352294 80058 352350
rect 79878 352170 79934 352226
rect 80002 352170 80058 352226
rect 79878 352046 79934 352102
rect 80002 352046 80058 352102
rect 79878 351922 79934 351978
rect 80002 351922 80058 351978
rect 78092 344402 78148 344458
rect 76524 307502 76580 307558
rect 83132 425402 83188 425458
rect 83132 404702 83188 404758
rect 80220 335762 80276 335818
rect 83132 374822 83188 374878
rect 79878 334294 79934 334350
rect 80002 334294 80058 334350
rect 79878 334170 79934 334226
rect 80002 334170 80058 334226
rect 79878 334046 79934 334102
rect 80002 334046 80058 334102
rect 79878 333922 79934 333978
rect 80002 333922 80058 333978
rect 79878 316294 79934 316350
rect 80002 316294 80058 316350
rect 79878 316170 79934 316226
rect 80002 316170 80058 316226
rect 79878 316046 79934 316102
rect 80002 316046 80058 316102
rect 79878 315922 79934 315978
rect 80002 315922 80058 315978
rect 79878 298294 79934 298350
rect 80002 298294 80058 298350
rect 79878 298170 79934 298226
rect 80002 298170 80058 298226
rect 79878 298046 79934 298102
rect 80002 298046 80058 298102
rect 79878 297922 79934 297978
rect 80002 297922 80058 297978
rect 78092 286802 78148 286858
rect 76524 285542 76580 285598
rect 70674 244294 70730 244350
rect 70798 244294 70854 244350
rect 70922 244294 70978 244350
rect 71046 244294 71102 244350
rect 70674 244170 70730 244226
rect 70798 244170 70854 244226
rect 70922 244170 70978 244226
rect 71046 244170 71102 244226
rect 70674 244046 70730 244102
rect 70798 244046 70854 244102
rect 70922 244046 70978 244102
rect 71046 244046 71102 244102
rect 70674 243922 70730 243978
rect 70798 243922 70854 243978
rect 70922 243922 70978 243978
rect 71046 243922 71102 243978
rect 66954 220294 67010 220350
rect 67078 220294 67134 220350
rect 67202 220294 67258 220350
rect 67326 220294 67382 220350
rect 66954 220170 67010 220226
rect 67078 220170 67134 220226
rect 67202 220170 67258 220226
rect 67326 220170 67382 220226
rect 66954 220046 67010 220102
rect 67078 220046 67134 220102
rect 67202 220046 67258 220102
rect 67326 220046 67382 220102
rect 66954 219922 67010 219978
rect 67078 219922 67134 219978
rect 67202 219922 67258 219978
rect 67326 219922 67382 219978
rect 64518 202294 64574 202350
rect 64642 202294 64698 202350
rect 64518 202170 64574 202226
rect 64642 202170 64698 202226
rect 64518 202046 64574 202102
rect 64642 202046 64698 202102
rect 64518 201922 64574 201978
rect 64642 201922 64698 201978
rect 66954 202294 67010 202350
rect 67078 202294 67134 202350
rect 67202 202294 67258 202350
rect 67326 202294 67382 202350
rect 66954 202170 67010 202226
rect 67078 202170 67134 202226
rect 67202 202170 67258 202226
rect 67326 202170 67382 202226
rect 66954 202046 67010 202102
rect 67078 202046 67134 202102
rect 67202 202046 67258 202102
rect 67326 202046 67382 202102
rect 66954 201922 67010 201978
rect 67078 201922 67134 201978
rect 67202 201922 67258 201978
rect 67326 201922 67382 201978
rect 62188 142622 62244 142678
rect 64518 184294 64574 184350
rect 64642 184294 64698 184350
rect 64518 184170 64574 184226
rect 64642 184170 64698 184226
rect 64518 184046 64574 184102
rect 64642 184046 64698 184102
rect 64518 183922 64574 183978
rect 64642 183922 64698 183978
rect 66954 184294 67010 184350
rect 67078 184294 67134 184350
rect 67202 184294 67258 184350
rect 67326 184294 67382 184350
rect 66954 184170 67010 184226
rect 67078 184170 67134 184226
rect 67202 184170 67258 184226
rect 67326 184170 67382 184226
rect 66954 184046 67010 184102
rect 67078 184046 67134 184102
rect 67202 184046 67258 184102
rect 67326 184046 67382 184102
rect 66954 183922 67010 183978
rect 67078 183922 67134 183978
rect 67202 183922 67258 183978
rect 67326 183922 67382 183978
rect 64518 166294 64574 166350
rect 64642 166294 64698 166350
rect 64518 166170 64574 166226
rect 64642 166170 64698 166226
rect 64518 166046 64574 166102
rect 64642 166046 64698 166102
rect 64518 165922 64574 165978
rect 64642 165922 64698 165978
rect 66954 166294 67010 166350
rect 67078 166294 67134 166350
rect 67202 166294 67258 166350
rect 67326 166294 67382 166350
rect 66954 166170 67010 166226
rect 67078 166170 67134 166226
rect 67202 166170 67258 166226
rect 67326 166170 67382 166226
rect 66954 166046 67010 166102
rect 67078 166046 67134 166102
rect 67202 166046 67258 166102
rect 67326 166046 67382 166102
rect 66954 165922 67010 165978
rect 67078 165922 67134 165978
rect 67202 165922 67258 165978
rect 67326 165922 67382 165978
rect 62748 142622 62804 142678
rect 66954 148294 67010 148350
rect 67078 148294 67134 148350
rect 67202 148294 67258 148350
rect 67326 148294 67382 148350
rect 66954 148170 67010 148226
rect 67078 148170 67134 148226
rect 67202 148170 67258 148226
rect 67326 148170 67382 148226
rect 66954 148046 67010 148102
rect 67078 148046 67134 148102
rect 67202 148046 67258 148102
rect 67326 148046 67382 148102
rect 66954 147922 67010 147978
rect 67078 147922 67134 147978
rect 67202 147922 67258 147978
rect 67326 147922 67382 147978
rect 63756 142262 63812 142318
rect 39954 136294 40010 136350
rect 40078 136294 40134 136350
rect 40202 136294 40258 136350
rect 40326 136294 40382 136350
rect 39954 136170 40010 136226
rect 40078 136170 40134 136226
rect 40202 136170 40258 136226
rect 40326 136170 40382 136226
rect 39954 136046 40010 136102
rect 40078 136046 40134 136102
rect 40202 136046 40258 136102
rect 40326 136046 40382 136102
rect 39954 135922 40010 135978
rect 40078 135922 40134 135978
rect 40202 135922 40258 135978
rect 40326 135922 40382 135978
rect 61130 130294 61186 130350
rect 61254 130294 61310 130350
rect 61378 130294 61434 130350
rect 61502 130294 61558 130350
rect 61130 130170 61186 130226
rect 61254 130170 61310 130226
rect 61378 130170 61434 130226
rect 61502 130170 61558 130226
rect 61130 130046 61186 130102
rect 61254 130046 61310 130102
rect 61378 130046 61434 130102
rect 61502 130046 61558 130102
rect 61130 129922 61186 129978
rect 61254 129922 61310 129978
rect 61378 129922 61434 129978
rect 61502 129922 61558 129978
rect 66954 130294 67010 130350
rect 67078 130294 67134 130350
rect 67202 130294 67258 130350
rect 67326 130294 67382 130350
rect 66954 130170 67010 130226
rect 67078 130170 67134 130226
rect 67202 130170 67258 130226
rect 67326 130170 67382 130226
rect 66954 130046 67010 130102
rect 67078 130046 67134 130102
rect 67202 130046 67258 130102
rect 67326 130046 67382 130102
rect 66954 129922 67010 129978
rect 67078 129922 67134 129978
rect 67202 129922 67258 129978
rect 67326 129922 67382 129978
rect 39954 118294 40010 118350
rect 40078 118294 40134 118350
rect 40202 118294 40258 118350
rect 40326 118294 40382 118350
rect 39954 118170 40010 118226
rect 40078 118170 40134 118226
rect 40202 118170 40258 118226
rect 40326 118170 40382 118226
rect 39954 118046 40010 118102
rect 40078 118046 40134 118102
rect 40202 118046 40258 118102
rect 40326 118046 40382 118102
rect 39954 117922 40010 117978
rect 40078 117922 40134 117978
rect 40202 117922 40258 117978
rect 40326 117922 40382 117978
rect 61930 118294 61986 118350
rect 62054 118294 62110 118350
rect 62178 118294 62234 118350
rect 62302 118294 62358 118350
rect 61930 118170 61986 118226
rect 62054 118170 62110 118226
rect 62178 118170 62234 118226
rect 62302 118170 62358 118226
rect 61930 118046 61986 118102
rect 62054 118046 62110 118102
rect 62178 118046 62234 118102
rect 62302 118046 62358 118102
rect 61930 117922 61986 117978
rect 62054 117922 62110 117978
rect 62178 117922 62234 117978
rect 62302 117922 62358 117978
rect 61130 112294 61186 112350
rect 61254 112294 61310 112350
rect 61378 112294 61434 112350
rect 61502 112294 61558 112350
rect 61130 112170 61186 112226
rect 61254 112170 61310 112226
rect 61378 112170 61434 112226
rect 61502 112170 61558 112226
rect 61130 112046 61186 112102
rect 61254 112046 61310 112102
rect 61378 112046 61434 112102
rect 61502 112046 61558 112102
rect 61130 111922 61186 111978
rect 61254 111922 61310 111978
rect 61378 111922 61434 111978
rect 61502 111922 61558 111978
rect 66954 112294 67010 112350
rect 67078 112294 67134 112350
rect 67202 112294 67258 112350
rect 67326 112294 67382 112350
rect 66954 112170 67010 112226
rect 67078 112170 67134 112226
rect 67202 112170 67258 112226
rect 67326 112170 67382 112226
rect 66954 112046 67010 112102
rect 67078 112046 67134 112102
rect 67202 112046 67258 112102
rect 67326 112046 67382 112102
rect 66954 111922 67010 111978
rect 67078 111922 67134 111978
rect 67202 111922 67258 111978
rect 67326 111922 67382 111978
rect 39954 100294 40010 100350
rect 40078 100294 40134 100350
rect 40202 100294 40258 100350
rect 40326 100294 40382 100350
rect 39954 100170 40010 100226
rect 40078 100170 40134 100226
rect 40202 100170 40258 100226
rect 40326 100170 40382 100226
rect 39954 100046 40010 100102
rect 40078 100046 40134 100102
rect 40202 100046 40258 100102
rect 40326 100046 40382 100102
rect 39954 99922 40010 99978
rect 40078 99922 40134 99978
rect 40202 99922 40258 99978
rect 40326 99922 40382 99978
rect 61930 100294 61986 100350
rect 62054 100294 62110 100350
rect 62178 100294 62234 100350
rect 62302 100294 62358 100350
rect 61930 100170 61986 100226
rect 62054 100170 62110 100226
rect 62178 100170 62234 100226
rect 62302 100170 62358 100226
rect 61930 100046 61986 100102
rect 62054 100046 62110 100102
rect 62178 100046 62234 100102
rect 62302 100046 62358 100102
rect 61930 99922 61986 99978
rect 62054 99922 62110 99978
rect 62178 99922 62234 99978
rect 62302 99922 62358 99978
rect 61130 94294 61186 94350
rect 61254 94294 61310 94350
rect 61378 94294 61434 94350
rect 61502 94294 61558 94350
rect 61130 94170 61186 94226
rect 61254 94170 61310 94226
rect 61378 94170 61434 94226
rect 61502 94170 61558 94226
rect 61130 94046 61186 94102
rect 61254 94046 61310 94102
rect 61378 94046 61434 94102
rect 61502 94046 61558 94102
rect 61130 93922 61186 93978
rect 61254 93922 61310 93978
rect 61378 93922 61434 93978
rect 61502 93922 61558 93978
rect 66954 94294 67010 94350
rect 67078 94294 67134 94350
rect 67202 94294 67258 94350
rect 67326 94294 67382 94350
rect 66954 94170 67010 94226
rect 67078 94170 67134 94226
rect 67202 94170 67258 94226
rect 67326 94170 67382 94226
rect 66954 94046 67010 94102
rect 67078 94046 67134 94102
rect 67202 94046 67258 94102
rect 67326 94046 67382 94102
rect 66954 93922 67010 93978
rect 67078 93922 67134 93978
rect 67202 93922 67258 93978
rect 67326 93922 67382 93978
rect 39954 82294 40010 82350
rect 40078 82294 40134 82350
rect 40202 82294 40258 82350
rect 40326 82294 40382 82350
rect 39954 82170 40010 82226
rect 40078 82170 40134 82226
rect 40202 82170 40258 82226
rect 40326 82170 40382 82226
rect 39954 82046 40010 82102
rect 40078 82046 40134 82102
rect 40202 82046 40258 82102
rect 40326 82046 40382 82102
rect 39954 81922 40010 81978
rect 40078 81922 40134 81978
rect 40202 81922 40258 81978
rect 40326 81922 40382 81978
rect 61930 82294 61986 82350
rect 62054 82294 62110 82350
rect 62178 82294 62234 82350
rect 62302 82294 62358 82350
rect 61930 82170 61986 82226
rect 62054 82170 62110 82226
rect 62178 82170 62234 82226
rect 62302 82170 62358 82226
rect 61930 82046 61986 82102
rect 62054 82046 62110 82102
rect 62178 82046 62234 82102
rect 62302 82046 62358 82102
rect 61930 81922 61986 81978
rect 62054 81922 62110 81978
rect 62178 81922 62234 81978
rect 62302 81922 62358 81978
rect 61130 76294 61186 76350
rect 61254 76294 61310 76350
rect 61378 76294 61434 76350
rect 61502 76294 61558 76350
rect 61130 76170 61186 76226
rect 61254 76170 61310 76226
rect 61378 76170 61434 76226
rect 61502 76170 61558 76226
rect 61130 76046 61186 76102
rect 61254 76046 61310 76102
rect 61378 76046 61434 76102
rect 61502 76046 61558 76102
rect 61130 75922 61186 75978
rect 61254 75922 61310 75978
rect 61378 75922 61434 75978
rect 61502 75922 61558 75978
rect 66954 76294 67010 76350
rect 67078 76294 67134 76350
rect 67202 76294 67258 76350
rect 67326 76294 67382 76350
rect 66954 76170 67010 76226
rect 67078 76170 67134 76226
rect 67202 76170 67258 76226
rect 67326 76170 67382 76226
rect 66954 76046 67010 76102
rect 67078 76046 67134 76102
rect 67202 76046 67258 76102
rect 67326 76046 67382 76102
rect 66954 75922 67010 75978
rect 67078 75922 67134 75978
rect 67202 75922 67258 75978
rect 67326 75922 67382 75978
rect 39954 64294 40010 64350
rect 40078 64294 40134 64350
rect 40202 64294 40258 64350
rect 40326 64294 40382 64350
rect 39954 64170 40010 64226
rect 40078 64170 40134 64226
rect 40202 64170 40258 64226
rect 40326 64170 40382 64226
rect 39954 64046 40010 64102
rect 40078 64046 40134 64102
rect 40202 64046 40258 64102
rect 40326 64046 40382 64102
rect 39954 63922 40010 63978
rect 40078 63922 40134 63978
rect 40202 63922 40258 63978
rect 40326 63922 40382 63978
rect 61930 64294 61986 64350
rect 62054 64294 62110 64350
rect 62178 64294 62234 64350
rect 62302 64294 62358 64350
rect 61930 64170 61986 64226
rect 62054 64170 62110 64226
rect 62178 64170 62234 64226
rect 62302 64170 62358 64226
rect 61930 64046 61986 64102
rect 62054 64046 62110 64102
rect 62178 64046 62234 64102
rect 62302 64046 62358 64102
rect 61930 63922 61986 63978
rect 62054 63922 62110 63978
rect 62178 63922 62234 63978
rect 62302 63922 62358 63978
rect 61130 58294 61186 58350
rect 61254 58294 61310 58350
rect 61378 58294 61434 58350
rect 61502 58294 61558 58350
rect 61130 58170 61186 58226
rect 61254 58170 61310 58226
rect 61378 58170 61434 58226
rect 61502 58170 61558 58226
rect 61130 58046 61186 58102
rect 61254 58046 61310 58102
rect 61378 58046 61434 58102
rect 61502 58046 61558 58102
rect 61130 57922 61186 57978
rect 61254 57922 61310 57978
rect 61378 57922 61434 57978
rect 61502 57922 61558 57978
rect 66954 58294 67010 58350
rect 67078 58294 67134 58350
rect 67202 58294 67258 58350
rect 67326 58294 67382 58350
rect 66954 58170 67010 58226
rect 67078 58170 67134 58226
rect 67202 58170 67258 58226
rect 67326 58170 67382 58226
rect 66954 58046 67010 58102
rect 67078 58046 67134 58102
rect 67202 58046 67258 58102
rect 67326 58046 67382 58102
rect 66954 57922 67010 57978
rect 67078 57922 67134 57978
rect 67202 57922 67258 57978
rect 67326 57922 67382 57978
rect 39954 46294 40010 46350
rect 40078 46294 40134 46350
rect 40202 46294 40258 46350
rect 40326 46294 40382 46350
rect 39954 46170 40010 46226
rect 40078 46170 40134 46226
rect 40202 46170 40258 46226
rect 40326 46170 40382 46226
rect 39954 46046 40010 46102
rect 40078 46046 40134 46102
rect 40202 46046 40258 46102
rect 40326 46046 40382 46102
rect 39954 45922 40010 45978
rect 40078 45922 40134 45978
rect 40202 45922 40258 45978
rect 40326 45922 40382 45978
rect 61930 46294 61986 46350
rect 62054 46294 62110 46350
rect 62178 46294 62234 46350
rect 62302 46294 62358 46350
rect 61930 46170 61986 46226
rect 62054 46170 62110 46226
rect 62178 46170 62234 46226
rect 62302 46170 62358 46226
rect 61930 46046 61986 46102
rect 62054 46046 62110 46102
rect 62178 46046 62234 46102
rect 62302 46046 62358 46102
rect 61930 45922 61986 45978
rect 62054 45922 62110 45978
rect 62178 45922 62234 45978
rect 62302 45922 62358 45978
rect 39954 28294 40010 28350
rect 40078 28294 40134 28350
rect 40202 28294 40258 28350
rect 40326 28294 40382 28350
rect 39954 28170 40010 28226
rect 40078 28170 40134 28226
rect 40202 28170 40258 28226
rect 40326 28170 40382 28226
rect 39954 28046 40010 28102
rect 40078 28046 40134 28102
rect 40202 28046 40258 28102
rect 40326 28046 40382 28102
rect 39954 27922 40010 27978
rect 40078 27922 40134 27978
rect 40202 27922 40258 27978
rect 40326 27922 40382 27978
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 66954 40294 67010 40350
rect 67078 40294 67134 40350
rect 67202 40294 67258 40350
rect 67326 40294 67382 40350
rect 66954 40170 67010 40226
rect 67078 40170 67134 40226
rect 67202 40170 67258 40226
rect 67326 40170 67382 40226
rect 66954 40046 67010 40102
rect 67078 40046 67134 40102
rect 67202 40046 67258 40102
rect 67326 40046 67382 40102
rect 66954 39922 67010 39978
rect 67078 39922 67134 39978
rect 67202 39922 67258 39978
rect 67326 39922 67382 39978
rect 66954 22294 67010 22350
rect 67078 22294 67134 22350
rect 67202 22294 67258 22350
rect 67326 22294 67382 22350
rect 66954 22170 67010 22226
rect 67078 22170 67134 22226
rect 67202 22170 67258 22226
rect 67326 22170 67382 22226
rect 66954 22046 67010 22102
rect 67078 22046 67134 22102
rect 67202 22046 67258 22102
rect 67326 22046 67382 22102
rect 66954 21922 67010 21978
rect 67078 21922 67134 21978
rect 67202 21922 67258 21978
rect 67326 21922 67382 21978
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 70674 226294 70730 226350
rect 70798 226294 70854 226350
rect 70922 226294 70978 226350
rect 71046 226294 71102 226350
rect 70674 226170 70730 226226
rect 70798 226170 70854 226226
rect 70922 226170 70978 226226
rect 71046 226170 71102 226226
rect 70674 226046 70730 226102
rect 70798 226046 70854 226102
rect 70922 226046 70978 226102
rect 71046 226046 71102 226102
rect 70674 225922 70730 225978
rect 70798 225922 70854 225978
rect 70922 225922 70978 225978
rect 71046 225922 71102 225978
rect 70674 208294 70730 208350
rect 70798 208294 70854 208350
rect 70922 208294 70978 208350
rect 71046 208294 71102 208350
rect 70674 208170 70730 208226
rect 70798 208170 70854 208226
rect 70922 208170 70978 208226
rect 71046 208170 71102 208226
rect 70674 208046 70730 208102
rect 70798 208046 70854 208102
rect 70922 208046 70978 208102
rect 71046 208046 71102 208102
rect 70674 207922 70730 207978
rect 70798 207922 70854 207978
rect 70922 207922 70978 207978
rect 71046 207922 71102 207978
rect 70674 190294 70730 190350
rect 70798 190294 70854 190350
rect 70922 190294 70978 190350
rect 71046 190294 71102 190350
rect 70674 190170 70730 190226
rect 70798 190170 70854 190226
rect 70922 190170 70978 190226
rect 71046 190170 71102 190226
rect 70674 190046 70730 190102
rect 70798 190046 70854 190102
rect 70922 190046 70978 190102
rect 71046 190046 71102 190102
rect 70674 189922 70730 189978
rect 70798 189922 70854 189978
rect 70922 189922 70978 189978
rect 71046 189922 71102 189978
rect 79878 190294 79934 190350
rect 80002 190294 80058 190350
rect 79878 190170 79934 190226
rect 80002 190170 80058 190226
rect 79878 190046 79934 190102
rect 80002 190046 80058 190102
rect 79878 189922 79934 189978
rect 80002 189922 80058 189978
rect 70674 172294 70730 172350
rect 70798 172294 70854 172350
rect 70922 172294 70978 172350
rect 71046 172294 71102 172350
rect 70674 172170 70730 172226
rect 70798 172170 70854 172226
rect 70922 172170 70978 172226
rect 71046 172170 71102 172226
rect 70674 172046 70730 172102
rect 70798 172046 70854 172102
rect 70922 172046 70978 172102
rect 71046 172046 71102 172102
rect 70674 171922 70730 171978
rect 70798 171922 70854 171978
rect 70922 171922 70978 171978
rect 71046 171922 71102 171978
rect 79878 172294 79934 172350
rect 80002 172294 80058 172350
rect 79878 172170 79934 172226
rect 80002 172170 80058 172226
rect 79878 172046 79934 172102
rect 80002 172046 80058 172102
rect 79878 171922 79934 171978
rect 80002 171922 80058 171978
rect 70674 154294 70730 154350
rect 70798 154294 70854 154350
rect 70922 154294 70978 154350
rect 71046 154294 71102 154350
rect 70674 154170 70730 154226
rect 70798 154170 70854 154226
rect 70922 154170 70978 154226
rect 71046 154170 71102 154226
rect 70674 154046 70730 154102
rect 70798 154046 70854 154102
rect 70922 154046 70978 154102
rect 71046 154046 71102 154102
rect 70674 153922 70730 153978
rect 70798 153922 70854 153978
rect 70922 153922 70978 153978
rect 71046 153922 71102 153978
rect 70674 136294 70730 136350
rect 70798 136294 70854 136350
rect 70922 136294 70978 136350
rect 71046 136294 71102 136350
rect 70674 136170 70730 136226
rect 70798 136170 70854 136226
rect 70922 136170 70978 136226
rect 71046 136170 71102 136226
rect 70674 136046 70730 136102
rect 70798 136046 70854 136102
rect 70922 136046 70978 136102
rect 71046 136046 71102 136102
rect 70674 135922 70730 135978
rect 70798 135922 70854 135978
rect 70922 135922 70978 135978
rect 71046 135922 71102 135978
rect 70674 118294 70730 118350
rect 70798 118294 70854 118350
rect 70922 118294 70978 118350
rect 71046 118294 71102 118350
rect 70674 118170 70730 118226
rect 70798 118170 70854 118226
rect 70922 118170 70978 118226
rect 71046 118170 71102 118226
rect 70674 118046 70730 118102
rect 70798 118046 70854 118102
rect 70922 118046 70978 118102
rect 71046 118046 71102 118102
rect 70674 117922 70730 117978
rect 70798 117922 70854 117978
rect 70922 117922 70978 117978
rect 71046 117922 71102 117978
rect 70674 100294 70730 100350
rect 70798 100294 70854 100350
rect 70922 100294 70978 100350
rect 71046 100294 71102 100350
rect 70674 100170 70730 100226
rect 70798 100170 70854 100226
rect 70922 100170 70978 100226
rect 71046 100170 71102 100226
rect 70674 100046 70730 100102
rect 70798 100046 70854 100102
rect 70922 100046 70978 100102
rect 71046 100046 71102 100102
rect 70674 99922 70730 99978
rect 70798 99922 70854 99978
rect 70922 99922 70978 99978
rect 71046 99922 71102 99978
rect 70674 82294 70730 82350
rect 70798 82294 70854 82350
rect 70922 82294 70978 82350
rect 71046 82294 71102 82350
rect 70674 82170 70730 82226
rect 70798 82170 70854 82226
rect 70922 82170 70978 82226
rect 71046 82170 71102 82226
rect 70674 82046 70730 82102
rect 70798 82046 70854 82102
rect 70922 82046 70978 82102
rect 71046 82046 71102 82102
rect 70674 81922 70730 81978
rect 70798 81922 70854 81978
rect 70922 81922 70978 81978
rect 71046 81922 71102 81978
rect 70674 64294 70730 64350
rect 70798 64294 70854 64350
rect 70922 64294 70978 64350
rect 71046 64294 71102 64350
rect 70674 64170 70730 64226
rect 70798 64170 70854 64226
rect 70922 64170 70978 64226
rect 71046 64170 71102 64226
rect 70674 64046 70730 64102
rect 70798 64046 70854 64102
rect 70922 64046 70978 64102
rect 71046 64046 71102 64102
rect 70674 63922 70730 63978
rect 70798 63922 70854 63978
rect 70922 63922 70978 63978
rect 71046 63922 71102 63978
rect 70674 46294 70730 46350
rect 70798 46294 70854 46350
rect 70922 46294 70978 46350
rect 71046 46294 71102 46350
rect 70674 46170 70730 46226
rect 70798 46170 70854 46226
rect 70922 46170 70978 46226
rect 71046 46170 71102 46226
rect 70674 46046 70730 46102
rect 70798 46046 70854 46102
rect 70922 46046 70978 46102
rect 71046 46046 71102 46102
rect 70674 45922 70730 45978
rect 70798 45922 70854 45978
rect 70922 45922 70978 45978
rect 71046 45922 71102 45978
rect 70674 28294 70730 28350
rect 70798 28294 70854 28350
rect 70922 28294 70978 28350
rect 71046 28294 71102 28350
rect 70674 28170 70730 28226
rect 70798 28170 70854 28226
rect 70922 28170 70978 28226
rect 71046 28170 71102 28226
rect 70674 28046 70730 28102
rect 70798 28046 70854 28102
rect 70922 28046 70978 28102
rect 71046 28046 71102 28102
rect 70674 27922 70730 27978
rect 70798 27922 70854 27978
rect 70922 27922 70978 27978
rect 71046 27922 71102 27978
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 83356 408122 83412 408178
rect 83468 425222 83524 425278
rect 83244 335942 83300 335998
rect 83356 374642 83412 374698
rect 101394 478294 101450 478350
rect 101518 478294 101574 478350
rect 101642 478294 101698 478350
rect 101766 478294 101822 478350
rect 101394 478170 101450 478226
rect 101518 478170 101574 478226
rect 101642 478170 101698 478226
rect 101766 478170 101822 478226
rect 101394 478046 101450 478102
rect 101518 478046 101574 478102
rect 101642 478046 101698 478102
rect 101766 478046 101822 478102
rect 101394 477922 101450 477978
rect 101518 477922 101574 477978
rect 101642 477922 101698 477978
rect 101766 477922 101822 477978
rect 101394 460294 101450 460350
rect 101518 460294 101574 460350
rect 101642 460294 101698 460350
rect 101766 460294 101822 460350
rect 101394 460170 101450 460226
rect 101518 460170 101574 460226
rect 101642 460170 101698 460226
rect 101766 460170 101822 460226
rect 101394 460046 101450 460102
rect 101518 460046 101574 460102
rect 101642 460046 101698 460102
rect 101766 460046 101822 460102
rect 101394 459922 101450 459978
rect 101518 459922 101574 459978
rect 101642 459922 101698 459978
rect 101766 459922 101822 459978
rect 101394 442294 101450 442350
rect 101518 442294 101574 442350
rect 101642 442294 101698 442350
rect 101766 442294 101822 442350
rect 101394 442170 101450 442226
rect 101518 442170 101574 442226
rect 101642 442170 101698 442226
rect 101766 442170 101822 442226
rect 101394 442046 101450 442102
rect 101518 442046 101574 442102
rect 101642 442046 101698 442102
rect 101766 442046 101822 442102
rect 101394 441922 101450 441978
rect 101518 441922 101574 441978
rect 101642 441922 101698 441978
rect 101766 441922 101822 441978
rect 128394 544294 128450 544350
rect 128518 544294 128574 544350
rect 128642 544294 128698 544350
rect 128766 544294 128822 544350
rect 128394 544170 128450 544226
rect 128518 544170 128574 544226
rect 128642 544170 128698 544226
rect 128766 544170 128822 544226
rect 128394 544046 128450 544102
rect 128518 544046 128574 544102
rect 128642 544046 128698 544102
rect 128766 544046 128822 544102
rect 128394 543922 128450 543978
rect 128518 543922 128574 543978
rect 128642 543922 128698 543978
rect 128766 543922 128822 543978
rect 128394 526294 128450 526350
rect 128518 526294 128574 526350
rect 128642 526294 128698 526350
rect 128766 526294 128822 526350
rect 128394 526170 128450 526226
rect 128518 526170 128574 526226
rect 128642 526170 128698 526226
rect 128766 526170 128822 526226
rect 128394 526046 128450 526102
rect 128518 526046 128574 526102
rect 128642 526046 128698 526102
rect 128766 526046 128822 526102
rect 128394 525922 128450 525978
rect 128518 525922 128574 525978
rect 128642 525922 128698 525978
rect 128766 525922 128822 525978
rect 128394 508294 128450 508350
rect 128518 508294 128574 508350
rect 128642 508294 128698 508350
rect 128766 508294 128822 508350
rect 128394 508170 128450 508226
rect 128518 508170 128574 508226
rect 128642 508170 128698 508226
rect 128766 508170 128822 508226
rect 128394 508046 128450 508102
rect 128518 508046 128574 508102
rect 128642 508046 128698 508102
rect 128766 508046 128822 508102
rect 128394 507922 128450 507978
rect 128518 507922 128574 507978
rect 128642 507922 128698 507978
rect 128766 507922 128822 507978
rect 128394 490294 128450 490350
rect 128518 490294 128574 490350
rect 128642 490294 128698 490350
rect 128766 490294 128822 490350
rect 128394 490170 128450 490226
rect 128518 490170 128574 490226
rect 128642 490170 128698 490226
rect 128766 490170 128822 490226
rect 128394 490046 128450 490102
rect 128518 490046 128574 490102
rect 128642 490046 128698 490102
rect 128766 490046 128822 490102
rect 128394 489922 128450 489978
rect 128518 489922 128574 489978
rect 128642 489922 128698 489978
rect 128766 489922 128822 489978
rect 128394 472294 128450 472350
rect 128518 472294 128574 472350
rect 128642 472294 128698 472350
rect 128766 472294 128822 472350
rect 128394 472170 128450 472226
rect 128518 472170 128574 472226
rect 128642 472170 128698 472226
rect 128766 472170 128822 472226
rect 128394 472046 128450 472102
rect 128518 472046 128574 472102
rect 128642 472046 128698 472102
rect 128766 472046 128822 472102
rect 128394 471922 128450 471978
rect 128518 471922 128574 471978
rect 128642 471922 128698 471978
rect 128766 471922 128822 471978
rect 128394 454294 128450 454350
rect 128518 454294 128574 454350
rect 128642 454294 128698 454350
rect 128766 454294 128822 454350
rect 128394 454170 128450 454226
rect 128518 454170 128574 454226
rect 128642 454170 128698 454226
rect 128766 454170 128822 454226
rect 128394 454046 128450 454102
rect 128518 454046 128574 454102
rect 128642 454046 128698 454102
rect 128766 454046 128822 454102
rect 128394 453922 128450 453978
rect 128518 453922 128574 453978
rect 128642 453922 128698 453978
rect 128766 453922 128822 453978
rect 128394 436294 128450 436350
rect 128518 436294 128574 436350
rect 128642 436294 128698 436350
rect 128766 436294 128822 436350
rect 128394 436170 128450 436226
rect 128518 436170 128574 436226
rect 128642 436170 128698 436226
rect 128766 436170 128822 436226
rect 128394 436046 128450 436102
rect 128518 436046 128574 436102
rect 128642 436046 128698 436102
rect 128766 436046 128822 436102
rect 128394 435922 128450 435978
rect 128518 435922 128574 435978
rect 128642 435922 128698 435978
rect 128766 435922 128822 435978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 132114 568294 132170 568350
rect 132238 568294 132294 568350
rect 132362 568294 132418 568350
rect 132486 568294 132542 568350
rect 132114 568170 132170 568226
rect 132238 568170 132294 568226
rect 132362 568170 132418 568226
rect 132486 568170 132542 568226
rect 132114 568046 132170 568102
rect 132238 568046 132294 568102
rect 132362 568046 132418 568102
rect 132486 568046 132542 568102
rect 132114 567922 132170 567978
rect 132238 567922 132294 567978
rect 132362 567922 132418 567978
rect 132486 567922 132542 567978
rect 132114 550294 132170 550350
rect 132238 550294 132294 550350
rect 132362 550294 132418 550350
rect 132486 550294 132542 550350
rect 132114 550170 132170 550226
rect 132238 550170 132294 550226
rect 132362 550170 132418 550226
rect 132486 550170 132542 550226
rect 132114 550046 132170 550102
rect 132238 550046 132294 550102
rect 132362 550046 132418 550102
rect 132486 550046 132542 550102
rect 132114 549922 132170 549978
rect 132238 549922 132294 549978
rect 132362 549922 132418 549978
rect 132486 549922 132542 549978
rect 132114 532294 132170 532350
rect 132238 532294 132294 532350
rect 132362 532294 132418 532350
rect 132486 532294 132542 532350
rect 132114 532170 132170 532226
rect 132238 532170 132294 532226
rect 132362 532170 132418 532226
rect 132486 532170 132542 532226
rect 132114 532046 132170 532102
rect 132238 532046 132294 532102
rect 132362 532046 132418 532102
rect 132486 532046 132542 532102
rect 132114 531922 132170 531978
rect 132238 531922 132294 531978
rect 132362 531922 132418 531978
rect 132486 531922 132542 531978
rect 132114 514294 132170 514350
rect 132238 514294 132294 514350
rect 132362 514294 132418 514350
rect 132486 514294 132542 514350
rect 132114 514170 132170 514226
rect 132238 514170 132294 514226
rect 132362 514170 132418 514226
rect 132486 514170 132542 514226
rect 132114 514046 132170 514102
rect 132238 514046 132294 514102
rect 132362 514046 132418 514102
rect 132486 514046 132542 514102
rect 132114 513922 132170 513978
rect 132238 513922 132294 513978
rect 132362 513922 132418 513978
rect 132486 513922 132542 513978
rect 132114 496294 132170 496350
rect 132238 496294 132294 496350
rect 132362 496294 132418 496350
rect 132486 496294 132542 496350
rect 132114 496170 132170 496226
rect 132238 496170 132294 496226
rect 132362 496170 132418 496226
rect 132486 496170 132542 496226
rect 132114 496046 132170 496102
rect 132238 496046 132294 496102
rect 132362 496046 132418 496102
rect 132486 496046 132542 496102
rect 132114 495922 132170 495978
rect 132238 495922 132294 495978
rect 132362 495922 132418 495978
rect 132486 495922 132542 495978
rect 132114 478294 132170 478350
rect 132238 478294 132294 478350
rect 132362 478294 132418 478350
rect 132486 478294 132542 478350
rect 132114 478170 132170 478226
rect 132238 478170 132294 478226
rect 132362 478170 132418 478226
rect 132486 478170 132542 478226
rect 132114 478046 132170 478102
rect 132238 478046 132294 478102
rect 132362 478046 132418 478102
rect 132486 478046 132542 478102
rect 132114 477922 132170 477978
rect 132238 477922 132294 477978
rect 132362 477922 132418 477978
rect 132486 477922 132542 477978
rect 132114 460294 132170 460350
rect 132238 460294 132294 460350
rect 132362 460294 132418 460350
rect 132486 460294 132542 460350
rect 132114 460170 132170 460226
rect 132238 460170 132294 460226
rect 132362 460170 132418 460226
rect 132486 460170 132542 460226
rect 132114 460046 132170 460102
rect 132238 460046 132294 460102
rect 132362 460046 132418 460102
rect 132486 460046 132542 460102
rect 132114 459922 132170 459978
rect 132238 459922 132294 459978
rect 132362 459922 132418 459978
rect 132486 459922 132542 459978
rect 132114 442294 132170 442350
rect 132238 442294 132294 442350
rect 132362 442294 132418 442350
rect 132486 442294 132542 442350
rect 132114 442170 132170 442226
rect 132238 442170 132294 442226
rect 132362 442170 132418 442226
rect 132486 442170 132542 442226
rect 132114 442046 132170 442102
rect 132238 442046 132294 442102
rect 132362 442046 132418 442102
rect 132486 442046 132542 442102
rect 132114 441922 132170 441978
rect 132238 441922 132294 441978
rect 132362 441922 132418 441978
rect 132486 441922 132542 441978
rect 159114 597156 159170 597212
rect 159238 597156 159294 597212
rect 159362 597156 159418 597212
rect 159486 597156 159542 597212
rect 159114 597032 159170 597088
rect 159238 597032 159294 597088
rect 159362 597032 159418 597088
rect 159486 597032 159542 597088
rect 159114 596908 159170 596964
rect 159238 596908 159294 596964
rect 159362 596908 159418 596964
rect 159486 596908 159542 596964
rect 159114 596784 159170 596840
rect 159238 596784 159294 596840
rect 159362 596784 159418 596840
rect 159486 596784 159542 596840
rect 159114 580294 159170 580350
rect 159238 580294 159294 580350
rect 159362 580294 159418 580350
rect 159486 580294 159542 580350
rect 159114 580170 159170 580226
rect 159238 580170 159294 580226
rect 159362 580170 159418 580226
rect 159486 580170 159542 580226
rect 159114 580046 159170 580102
rect 159238 580046 159294 580102
rect 159362 580046 159418 580102
rect 159486 580046 159542 580102
rect 159114 579922 159170 579978
rect 159238 579922 159294 579978
rect 159362 579922 159418 579978
rect 159486 579922 159542 579978
rect 159114 562294 159170 562350
rect 159238 562294 159294 562350
rect 159362 562294 159418 562350
rect 159486 562294 159542 562350
rect 159114 562170 159170 562226
rect 159238 562170 159294 562226
rect 159362 562170 159418 562226
rect 159486 562170 159542 562226
rect 159114 562046 159170 562102
rect 159238 562046 159294 562102
rect 159362 562046 159418 562102
rect 159486 562046 159542 562102
rect 159114 561922 159170 561978
rect 159238 561922 159294 561978
rect 159362 561922 159418 561978
rect 159486 561922 159542 561978
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 162834 568294 162890 568350
rect 162958 568294 163014 568350
rect 163082 568294 163138 568350
rect 163206 568294 163262 568350
rect 162834 568170 162890 568226
rect 162958 568170 163014 568226
rect 163082 568170 163138 568226
rect 163206 568170 163262 568226
rect 162834 568046 162890 568102
rect 162958 568046 163014 568102
rect 163082 568046 163138 568102
rect 163206 568046 163262 568102
rect 162834 567922 162890 567978
rect 162958 567922 163014 567978
rect 163082 567922 163138 567978
rect 163206 567922 163262 567978
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 189834 562294 189890 562350
rect 189958 562294 190014 562350
rect 190082 562294 190138 562350
rect 190206 562294 190262 562350
rect 189834 562170 189890 562226
rect 189958 562170 190014 562226
rect 190082 562170 190138 562226
rect 190206 562170 190262 562226
rect 189834 562046 189890 562102
rect 189958 562046 190014 562102
rect 190082 562046 190138 562102
rect 190206 562046 190262 562102
rect 189834 561922 189890 561978
rect 189958 561922 190014 561978
rect 190082 561922 190138 561978
rect 190206 561922 190262 561978
rect 162834 550294 162890 550350
rect 162958 550294 163014 550350
rect 163082 550294 163138 550350
rect 163206 550294 163262 550350
rect 162834 550170 162890 550226
rect 162958 550170 163014 550226
rect 163082 550170 163138 550226
rect 163206 550170 163262 550226
rect 162834 550046 162890 550102
rect 162958 550046 163014 550102
rect 163082 550046 163138 550102
rect 163206 550046 163262 550102
rect 162834 549922 162890 549978
rect 162958 549922 163014 549978
rect 163082 549922 163138 549978
rect 163206 549922 163262 549978
rect 179878 550294 179934 550350
rect 180002 550294 180058 550350
rect 179878 550170 179934 550226
rect 180002 550170 180058 550226
rect 179878 550046 179934 550102
rect 180002 550046 180058 550102
rect 179878 549922 179934 549978
rect 180002 549922 180058 549978
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 193554 568294 193610 568350
rect 193678 568294 193734 568350
rect 193802 568294 193858 568350
rect 193926 568294 193982 568350
rect 193554 568170 193610 568226
rect 193678 568170 193734 568226
rect 193802 568170 193858 568226
rect 193926 568170 193982 568226
rect 193554 568046 193610 568102
rect 193678 568046 193734 568102
rect 193802 568046 193858 568102
rect 193926 568046 193982 568102
rect 193554 567922 193610 567978
rect 193678 567922 193734 567978
rect 193802 567922 193858 567978
rect 193926 567922 193982 567978
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 220554 562294 220610 562350
rect 220678 562294 220734 562350
rect 220802 562294 220858 562350
rect 220926 562294 220982 562350
rect 220554 562170 220610 562226
rect 220678 562170 220734 562226
rect 220802 562170 220858 562226
rect 220926 562170 220982 562226
rect 220554 562046 220610 562102
rect 220678 562046 220734 562102
rect 220802 562046 220858 562102
rect 220926 562046 220982 562102
rect 220554 561922 220610 561978
rect 220678 561922 220734 561978
rect 220802 561922 220858 561978
rect 220926 561922 220982 561978
rect 193554 550294 193610 550350
rect 193678 550294 193734 550350
rect 193802 550294 193858 550350
rect 193926 550294 193982 550350
rect 193554 550170 193610 550226
rect 193678 550170 193734 550226
rect 193802 550170 193858 550226
rect 193926 550170 193982 550226
rect 193554 550046 193610 550102
rect 193678 550046 193734 550102
rect 193802 550046 193858 550102
rect 193926 550046 193982 550102
rect 193554 549922 193610 549978
rect 193678 549922 193734 549978
rect 193802 549922 193858 549978
rect 193926 549922 193982 549978
rect 210598 550294 210654 550350
rect 210722 550294 210778 550350
rect 210598 550170 210654 550226
rect 210722 550170 210778 550226
rect 210598 550046 210654 550102
rect 210722 550046 210778 550102
rect 210598 549922 210654 549978
rect 210722 549922 210778 549978
rect 159114 544294 159170 544350
rect 159238 544294 159294 544350
rect 159362 544294 159418 544350
rect 159486 544294 159542 544350
rect 159114 544170 159170 544226
rect 159238 544170 159294 544226
rect 159362 544170 159418 544226
rect 159486 544170 159542 544226
rect 159114 544046 159170 544102
rect 159238 544046 159294 544102
rect 159362 544046 159418 544102
rect 159486 544046 159542 544102
rect 159114 543922 159170 543978
rect 159238 543922 159294 543978
rect 159362 543922 159418 543978
rect 159486 543922 159542 543978
rect 164518 544294 164574 544350
rect 164642 544294 164698 544350
rect 164518 544170 164574 544226
rect 164642 544170 164698 544226
rect 164518 544046 164574 544102
rect 164642 544046 164698 544102
rect 164518 543922 164574 543978
rect 164642 543922 164698 543978
rect 195238 544294 195294 544350
rect 195362 544294 195418 544350
rect 195238 544170 195294 544226
rect 195362 544170 195418 544226
rect 195238 544046 195294 544102
rect 195362 544046 195418 544102
rect 195238 543922 195294 543978
rect 195362 543922 195418 543978
rect 179878 532294 179934 532350
rect 180002 532294 180058 532350
rect 179878 532170 179934 532226
rect 180002 532170 180058 532226
rect 179878 532046 179934 532102
rect 180002 532046 180058 532102
rect 179878 531922 179934 531978
rect 180002 531922 180058 531978
rect 210598 532294 210654 532350
rect 210722 532294 210778 532350
rect 210598 532170 210654 532226
rect 210722 532170 210778 532226
rect 210598 532046 210654 532102
rect 210722 532046 210778 532102
rect 210598 531922 210654 531978
rect 210722 531922 210778 531978
rect 159114 526294 159170 526350
rect 159238 526294 159294 526350
rect 159362 526294 159418 526350
rect 159486 526294 159542 526350
rect 159114 526170 159170 526226
rect 159238 526170 159294 526226
rect 159362 526170 159418 526226
rect 159486 526170 159542 526226
rect 159114 526046 159170 526102
rect 159238 526046 159294 526102
rect 159362 526046 159418 526102
rect 159486 526046 159542 526102
rect 159114 525922 159170 525978
rect 159238 525922 159294 525978
rect 159362 525922 159418 525978
rect 159486 525922 159542 525978
rect 164518 526294 164574 526350
rect 164642 526294 164698 526350
rect 164518 526170 164574 526226
rect 164642 526170 164698 526226
rect 164518 526046 164574 526102
rect 164642 526046 164698 526102
rect 164518 525922 164574 525978
rect 164642 525922 164698 525978
rect 195238 526294 195294 526350
rect 195362 526294 195418 526350
rect 195238 526170 195294 526226
rect 195362 526170 195418 526226
rect 195238 526046 195294 526102
rect 195362 526046 195418 526102
rect 195238 525922 195294 525978
rect 195362 525922 195418 525978
rect 179878 514294 179934 514350
rect 180002 514294 180058 514350
rect 179878 514170 179934 514226
rect 180002 514170 180058 514226
rect 179878 514046 179934 514102
rect 180002 514046 180058 514102
rect 179878 513922 179934 513978
rect 180002 513922 180058 513978
rect 210598 514294 210654 514350
rect 210722 514294 210778 514350
rect 210598 514170 210654 514226
rect 210722 514170 210778 514226
rect 210598 514046 210654 514102
rect 210722 514046 210778 514102
rect 210598 513922 210654 513978
rect 210722 513922 210778 513978
rect 159114 508294 159170 508350
rect 159238 508294 159294 508350
rect 159362 508294 159418 508350
rect 159486 508294 159542 508350
rect 159114 508170 159170 508226
rect 159238 508170 159294 508226
rect 159362 508170 159418 508226
rect 159486 508170 159542 508226
rect 159114 508046 159170 508102
rect 159238 508046 159294 508102
rect 159362 508046 159418 508102
rect 159486 508046 159542 508102
rect 159114 507922 159170 507978
rect 159238 507922 159294 507978
rect 159362 507922 159418 507978
rect 159486 507922 159542 507978
rect 164518 508294 164574 508350
rect 164642 508294 164698 508350
rect 164518 508170 164574 508226
rect 164642 508170 164698 508226
rect 164518 508046 164574 508102
rect 164642 508046 164698 508102
rect 164518 507922 164574 507978
rect 164642 507922 164698 507978
rect 195238 508294 195294 508350
rect 195362 508294 195418 508350
rect 195238 508170 195294 508226
rect 195362 508170 195418 508226
rect 195238 508046 195294 508102
rect 195362 508046 195418 508102
rect 195238 507922 195294 507978
rect 195362 507922 195418 507978
rect 159114 490294 159170 490350
rect 159238 490294 159294 490350
rect 159362 490294 159418 490350
rect 159486 490294 159542 490350
rect 159114 490170 159170 490226
rect 159238 490170 159294 490226
rect 159362 490170 159418 490226
rect 159486 490170 159542 490226
rect 159114 490046 159170 490102
rect 159238 490046 159294 490102
rect 159362 490046 159418 490102
rect 159486 490046 159542 490102
rect 159114 489922 159170 489978
rect 159238 489922 159294 489978
rect 159362 489922 159418 489978
rect 159486 489922 159542 489978
rect 159114 472294 159170 472350
rect 159238 472294 159294 472350
rect 159362 472294 159418 472350
rect 159486 472294 159542 472350
rect 159114 472170 159170 472226
rect 159238 472170 159294 472226
rect 159362 472170 159418 472226
rect 159486 472170 159542 472226
rect 159114 472046 159170 472102
rect 159238 472046 159294 472102
rect 159362 472046 159418 472102
rect 159486 472046 159542 472102
rect 159114 471922 159170 471978
rect 159238 471922 159294 471978
rect 159362 471922 159418 471978
rect 159486 471922 159542 471978
rect 159114 454294 159170 454350
rect 159238 454294 159294 454350
rect 159362 454294 159418 454350
rect 159486 454294 159542 454350
rect 159114 454170 159170 454226
rect 159238 454170 159294 454226
rect 159362 454170 159418 454226
rect 159486 454170 159542 454226
rect 159114 454046 159170 454102
rect 159238 454046 159294 454102
rect 159362 454046 159418 454102
rect 159486 454046 159542 454102
rect 159114 453922 159170 453978
rect 159238 453922 159294 453978
rect 159362 453922 159418 453978
rect 159486 453922 159542 453978
rect 159114 436294 159170 436350
rect 159238 436294 159294 436350
rect 159362 436294 159418 436350
rect 159486 436294 159542 436350
rect 159114 436170 159170 436226
rect 159238 436170 159294 436226
rect 159362 436170 159418 436226
rect 159486 436170 159542 436226
rect 159114 436046 159170 436102
rect 159238 436046 159294 436102
rect 159362 436046 159418 436102
rect 159486 436046 159542 436102
rect 159114 435922 159170 435978
rect 159238 435922 159294 435978
rect 159362 435922 159418 435978
rect 159486 435922 159542 435978
rect 162834 496294 162890 496350
rect 162958 496294 163014 496350
rect 163082 496294 163138 496350
rect 163206 496294 163262 496350
rect 162834 496170 162890 496226
rect 162958 496170 163014 496226
rect 163082 496170 163138 496226
rect 163206 496170 163262 496226
rect 162834 496046 162890 496102
rect 162958 496046 163014 496102
rect 163082 496046 163138 496102
rect 163206 496046 163262 496102
rect 162834 495922 162890 495978
rect 162958 495922 163014 495978
rect 163082 495922 163138 495978
rect 163206 495922 163262 495978
rect 189834 490294 189890 490350
rect 189958 490294 190014 490350
rect 190082 490294 190138 490350
rect 190206 490294 190262 490350
rect 189834 490170 189890 490226
rect 189958 490170 190014 490226
rect 190082 490170 190138 490226
rect 190206 490170 190262 490226
rect 189834 490046 189890 490102
rect 189958 490046 190014 490102
rect 190082 490046 190138 490102
rect 190206 490046 190262 490102
rect 189834 489922 189890 489978
rect 189958 489922 190014 489978
rect 190082 489922 190138 489978
rect 190206 489922 190262 489978
rect 169596 488042 169652 488098
rect 162834 478294 162890 478350
rect 162958 478294 163014 478350
rect 163082 478294 163138 478350
rect 163206 478294 163262 478350
rect 162834 478170 162890 478226
rect 162958 478170 163014 478226
rect 163082 478170 163138 478226
rect 163206 478170 163262 478226
rect 162834 478046 162890 478102
rect 162958 478046 163014 478102
rect 163082 478046 163138 478102
rect 163206 478046 163262 478102
rect 162834 477922 162890 477978
rect 162958 477922 163014 477978
rect 163082 477922 163138 477978
rect 163206 477922 163262 477978
rect 166236 479582 166292 479638
rect 162834 460294 162890 460350
rect 162958 460294 163014 460350
rect 163082 460294 163138 460350
rect 163206 460294 163262 460350
rect 162834 460170 162890 460226
rect 162958 460170 163014 460226
rect 163082 460170 163138 460226
rect 163206 460170 163262 460226
rect 162834 460046 162890 460102
rect 162958 460046 163014 460102
rect 163082 460046 163138 460102
rect 163206 460046 163262 460102
rect 162834 459922 162890 459978
rect 162958 459922 163014 459978
rect 163082 459922 163138 459978
rect 163206 459922 163262 459978
rect 162834 442294 162890 442350
rect 162958 442294 163014 442350
rect 163082 442294 163138 442350
rect 163206 442294 163262 442350
rect 162834 442170 162890 442226
rect 162958 442170 163014 442226
rect 163082 442170 163138 442226
rect 163206 442170 163262 442226
rect 162834 442046 162890 442102
rect 162958 442046 163014 442102
rect 163082 442046 163138 442102
rect 163206 442046 163262 442102
rect 162834 441922 162890 441978
rect 162958 441922 163014 441978
rect 163082 441922 163138 441978
rect 163206 441922 163262 441978
rect 164556 472562 164612 472618
rect 189834 472294 189890 472350
rect 189958 472294 190014 472350
rect 190082 472294 190138 472350
rect 190206 472294 190262 472350
rect 189834 472170 189890 472226
rect 189958 472170 190014 472226
rect 190082 472170 190138 472226
rect 190206 472170 190262 472226
rect 189834 472046 189890 472102
rect 189958 472046 190014 472102
rect 190082 472046 190138 472102
rect 190206 472046 190262 472102
rect 189834 471922 189890 471978
rect 189958 471922 190014 471978
rect 190082 471922 190138 471978
rect 190206 471922 190262 471978
rect 189834 454294 189890 454350
rect 189958 454294 190014 454350
rect 190082 454294 190138 454350
rect 190206 454294 190262 454350
rect 189834 454170 189890 454226
rect 189958 454170 190014 454226
rect 190082 454170 190138 454226
rect 190206 454170 190262 454226
rect 189834 454046 189890 454102
rect 189958 454046 190014 454102
rect 190082 454046 190138 454102
rect 190206 454046 190262 454102
rect 189834 453922 189890 453978
rect 189958 453922 190014 453978
rect 190082 453922 190138 453978
rect 190206 453922 190262 453978
rect 189834 436294 189890 436350
rect 189958 436294 190014 436350
rect 190082 436294 190138 436350
rect 190206 436294 190262 436350
rect 189834 436170 189890 436226
rect 189958 436170 190014 436226
rect 190082 436170 190138 436226
rect 190206 436170 190262 436226
rect 189834 436046 189890 436102
rect 189958 436046 190014 436102
rect 190082 436046 190138 436102
rect 190206 436046 190262 436102
rect 189834 435922 189890 435978
rect 189958 435922 190014 435978
rect 190082 435922 190138 435978
rect 190206 435922 190262 435978
rect 193554 496294 193610 496350
rect 193678 496294 193734 496350
rect 193802 496294 193858 496350
rect 193926 496294 193982 496350
rect 193554 496170 193610 496226
rect 193678 496170 193734 496226
rect 193802 496170 193858 496226
rect 193926 496170 193982 496226
rect 193554 496046 193610 496102
rect 193678 496046 193734 496102
rect 193802 496046 193858 496102
rect 193926 496046 193982 496102
rect 193554 495922 193610 495978
rect 193678 495922 193734 495978
rect 193802 495922 193858 495978
rect 193926 495922 193982 495978
rect 193554 478294 193610 478350
rect 193678 478294 193734 478350
rect 193802 478294 193858 478350
rect 193926 478294 193982 478350
rect 193554 478170 193610 478226
rect 193678 478170 193734 478226
rect 193802 478170 193858 478226
rect 193926 478170 193982 478226
rect 193554 478046 193610 478102
rect 193678 478046 193734 478102
rect 193802 478046 193858 478102
rect 193926 478046 193982 478102
rect 193554 477922 193610 477978
rect 193678 477922 193734 477978
rect 193802 477922 193858 477978
rect 193926 477922 193982 477978
rect 193554 460294 193610 460350
rect 193678 460294 193734 460350
rect 193802 460294 193858 460350
rect 193926 460294 193982 460350
rect 193554 460170 193610 460226
rect 193678 460170 193734 460226
rect 193802 460170 193858 460226
rect 193926 460170 193982 460226
rect 193554 460046 193610 460102
rect 193678 460046 193734 460102
rect 193802 460046 193858 460102
rect 193926 460046 193982 460102
rect 193554 459922 193610 459978
rect 193678 459922 193734 459978
rect 193802 459922 193858 459978
rect 193926 459922 193982 459978
rect 193554 442294 193610 442350
rect 193678 442294 193734 442350
rect 193802 442294 193858 442350
rect 193926 442294 193982 442350
rect 193554 442170 193610 442226
rect 193678 442170 193734 442226
rect 193802 442170 193858 442226
rect 193926 442170 193982 442226
rect 193554 442046 193610 442102
rect 193678 442046 193734 442102
rect 193802 442046 193858 442102
rect 193926 442046 193982 442102
rect 193554 441922 193610 441978
rect 193678 441922 193734 441978
rect 193802 441922 193858 441978
rect 193926 441922 193982 441978
rect 220554 544294 220610 544350
rect 220678 544294 220734 544350
rect 220802 544294 220858 544350
rect 220926 544294 220982 544350
rect 220554 544170 220610 544226
rect 220678 544170 220734 544226
rect 220802 544170 220858 544226
rect 220926 544170 220982 544226
rect 220554 544046 220610 544102
rect 220678 544046 220734 544102
rect 220802 544046 220858 544102
rect 220926 544046 220982 544102
rect 220554 543922 220610 543978
rect 220678 543922 220734 543978
rect 220802 543922 220858 543978
rect 220926 543922 220982 543978
rect 220554 526294 220610 526350
rect 220678 526294 220734 526350
rect 220802 526294 220858 526350
rect 220926 526294 220982 526350
rect 220554 526170 220610 526226
rect 220678 526170 220734 526226
rect 220802 526170 220858 526226
rect 220926 526170 220982 526226
rect 220554 526046 220610 526102
rect 220678 526046 220734 526102
rect 220802 526046 220858 526102
rect 220926 526046 220982 526102
rect 220554 525922 220610 525978
rect 220678 525922 220734 525978
rect 220802 525922 220858 525978
rect 220926 525922 220982 525978
rect 220554 508294 220610 508350
rect 220678 508294 220734 508350
rect 220802 508294 220858 508350
rect 220926 508294 220982 508350
rect 220554 508170 220610 508226
rect 220678 508170 220734 508226
rect 220802 508170 220858 508226
rect 220926 508170 220982 508226
rect 220554 508046 220610 508102
rect 220678 508046 220734 508102
rect 220802 508046 220858 508102
rect 220926 508046 220982 508102
rect 220554 507922 220610 507978
rect 220678 507922 220734 507978
rect 220802 507922 220858 507978
rect 220926 507922 220982 507978
rect 220554 490294 220610 490350
rect 220678 490294 220734 490350
rect 220802 490294 220858 490350
rect 220926 490294 220982 490350
rect 220554 490170 220610 490226
rect 220678 490170 220734 490226
rect 220802 490170 220858 490226
rect 220926 490170 220982 490226
rect 220554 490046 220610 490102
rect 220678 490046 220734 490102
rect 220802 490046 220858 490102
rect 220926 490046 220982 490102
rect 220554 489922 220610 489978
rect 220678 489922 220734 489978
rect 220802 489922 220858 489978
rect 220926 489922 220982 489978
rect 220554 472294 220610 472350
rect 220678 472294 220734 472350
rect 220802 472294 220858 472350
rect 220926 472294 220982 472350
rect 220554 472170 220610 472226
rect 220678 472170 220734 472226
rect 220802 472170 220858 472226
rect 220926 472170 220982 472226
rect 220554 472046 220610 472102
rect 220678 472046 220734 472102
rect 220802 472046 220858 472102
rect 220926 472046 220982 472102
rect 220554 471922 220610 471978
rect 220678 471922 220734 471978
rect 220802 471922 220858 471978
rect 220926 471922 220982 471978
rect 220554 454294 220610 454350
rect 220678 454294 220734 454350
rect 220802 454294 220858 454350
rect 220926 454294 220982 454350
rect 220554 454170 220610 454226
rect 220678 454170 220734 454226
rect 220802 454170 220858 454226
rect 220926 454170 220982 454226
rect 220554 454046 220610 454102
rect 220678 454046 220734 454102
rect 220802 454046 220858 454102
rect 220926 454046 220982 454102
rect 220554 453922 220610 453978
rect 220678 453922 220734 453978
rect 220802 453922 220858 453978
rect 220926 453922 220982 453978
rect 220554 436294 220610 436350
rect 220678 436294 220734 436350
rect 220802 436294 220858 436350
rect 220926 436294 220982 436350
rect 220554 436170 220610 436226
rect 220678 436170 220734 436226
rect 220802 436170 220858 436226
rect 220926 436170 220982 436226
rect 220554 436046 220610 436102
rect 220678 436046 220734 436102
rect 220802 436046 220858 436102
rect 220926 436046 220982 436102
rect 220554 435922 220610 435978
rect 220678 435922 220734 435978
rect 220802 435922 220858 435978
rect 220926 435922 220982 435978
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 224274 568294 224330 568350
rect 224398 568294 224454 568350
rect 224522 568294 224578 568350
rect 224646 568294 224702 568350
rect 224274 568170 224330 568226
rect 224398 568170 224454 568226
rect 224522 568170 224578 568226
rect 224646 568170 224702 568226
rect 224274 568046 224330 568102
rect 224398 568046 224454 568102
rect 224522 568046 224578 568102
rect 224646 568046 224702 568102
rect 224274 567922 224330 567978
rect 224398 567922 224454 567978
rect 224522 567922 224578 567978
rect 224646 567922 224702 567978
rect 224274 550294 224330 550350
rect 224398 550294 224454 550350
rect 224522 550294 224578 550350
rect 224646 550294 224702 550350
rect 224274 550170 224330 550226
rect 224398 550170 224454 550226
rect 224522 550170 224578 550226
rect 224646 550170 224702 550226
rect 224274 550046 224330 550102
rect 224398 550046 224454 550102
rect 224522 550046 224578 550102
rect 224646 550046 224702 550102
rect 224274 549922 224330 549978
rect 224398 549922 224454 549978
rect 224522 549922 224578 549978
rect 224646 549922 224702 549978
rect 224274 532294 224330 532350
rect 224398 532294 224454 532350
rect 224522 532294 224578 532350
rect 224646 532294 224702 532350
rect 224274 532170 224330 532226
rect 224398 532170 224454 532226
rect 224522 532170 224578 532226
rect 224646 532170 224702 532226
rect 224274 532046 224330 532102
rect 224398 532046 224454 532102
rect 224522 532046 224578 532102
rect 224646 532046 224702 532102
rect 224274 531922 224330 531978
rect 224398 531922 224454 531978
rect 224522 531922 224578 531978
rect 224646 531922 224702 531978
rect 224274 514294 224330 514350
rect 224398 514294 224454 514350
rect 224522 514294 224578 514350
rect 224646 514294 224702 514350
rect 224274 514170 224330 514226
rect 224398 514170 224454 514226
rect 224522 514170 224578 514226
rect 224646 514170 224702 514226
rect 224274 514046 224330 514102
rect 224398 514046 224454 514102
rect 224522 514046 224578 514102
rect 224646 514046 224702 514102
rect 224274 513922 224330 513978
rect 224398 513922 224454 513978
rect 224522 513922 224578 513978
rect 224646 513922 224702 513978
rect 224274 496294 224330 496350
rect 224398 496294 224454 496350
rect 224522 496294 224578 496350
rect 224646 496294 224702 496350
rect 224274 496170 224330 496226
rect 224398 496170 224454 496226
rect 224522 496170 224578 496226
rect 224646 496170 224702 496226
rect 224274 496046 224330 496102
rect 224398 496046 224454 496102
rect 224522 496046 224578 496102
rect 224646 496046 224702 496102
rect 224274 495922 224330 495978
rect 224398 495922 224454 495978
rect 224522 495922 224578 495978
rect 224646 495922 224702 495978
rect 224274 478294 224330 478350
rect 224398 478294 224454 478350
rect 224522 478294 224578 478350
rect 224646 478294 224702 478350
rect 224274 478170 224330 478226
rect 224398 478170 224454 478226
rect 224522 478170 224578 478226
rect 224646 478170 224702 478226
rect 224274 478046 224330 478102
rect 224398 478046 224454 478102
rect 224522 478046 224578 478102
rect 224646 478046 224702 478102
rect 224274 477922 224330 477978
rect 224398 477922 224454 477978
rect 224522 477922 224578 477978
rect 224646 477922 224702 477978
rect 224274 460294 224330 460350
rect 224398 460294 224454 460350
rect 224522 460294 224578 460350
rect 224646 460294 224702 460350
rect 224274 460170 224330 460226
rect 224398 460170 224454 460226
rect 224522 460170 224578 460226
rect 224646 460170 224702 460226
rect 224274 460046 224330 460102
rect 224398 460046 224454 460102
rect 224522 460046 224578 460102
rect 224646 460046 224702 460102
rect 224274 459922 224330 459978
rect 224398 459922 224454 459978
rect 224522 459922 224578 459978
rect 224646 459922 224702 459978
rect 224274 442294 224330 442350
rect 224398 442294 224454 442350
rect 224522 442294 224578 442350
rect 224646 442294 224702 442350
rect 224274 442170 224330 442226
rect 224398 442170 224454 442226
rect 224522 442170 224578 442226
rect 224646 442170 224702 442226
rect 224274 442046 224330 442102
rect 224398 442046 224454 442102
rect 224522 442046 224578 442102
rect 224646 442046 224702 442102
rect 224274 441922 224330 441978
rect 224398 441922 224454 441978
rect 224522 441922 224578 441978
rect 224646 441922 224702 441978
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 251274 562294 251330 562350
rect 251398 562294 251454 562350
rect 251522 562294 251578 562350
rect 251646 562294 251702 562350
rect 251274 562170 251330 562226
rect 251398 562170 251454 562226
rect 251522 562170 251578 562226
rect 251646 562170 251702 562226
rect 251274 562046 251330 562102
rect 251398 562046 251454 562102
rect 251522 562046 251578 562102
rect 251646 562046 251702 562102
rect 251274 561922 251330 561978
rect 251398 561922 251454 561978
rect 251522 561922 251578 561978
rect 251646 561922 251702 561978
rect 251274 544294 251330 544350
rect 251398 544294 251454 544350
rect 251522 544294 251578 544350
rect 251646 544294 251702 544350
rect 251274 544170 251330 544226
rect 251398 544170 251454 544226
rect 251522 544170 251578 544226
rect 251646 544170 251702 544226
rect 251274 544046 251330 544102
rect 251398 544046 251454 544102
rect 251522 544046 251578 544102
rect 251646 544046 251702 544102
rect 251274 543922 251330 543978
rect 251398 543922 251454 543978
rect 251522 543922 251578 543978
rect 251646 543922 251702 543978
rect 251274 526294 251330 526350
rect 251398 526294 251454 526350
rect 251522 526294 251578 526350
rect 251646 526294 251702 526350
rect 251274 526170 251330 526226
rect 251398 526170 251454 526226
rect 251522 526170 251578 526226
rect 251646 526170 251702 526226
rect 251274 526046 251330 526102
rect 251398 526046 251454 526102
rect 251522 526046 251578 526102
rect 251646 526046 251702 526102
rect 251274 525922 251330 525978
rect 251398 525922 251454 525978
rect 251522 525922 251578 525978
rect 251646 525922 251702 525978
rect 251274 508294 251330 508350
rect 251398 508294 251454 508350
rect 251522 508294 251578 508350
rect 251646 508294 251702 508350
rect 251274 508170 251330 508226
rect 251398 508170 251454 508226
rect 251522 508170 251578 508226
rect 251646 508170 251702 508226
rect 251274 508046 251330 508102
rect 251398 508046 251454 508102
rect 251522 508046 251578 508102
rect 251646 508046 251702 508102
rect 251274 507922 251330 507978
rect 251398 507922 251454 507978
rect 251522 507922 251578 507978
rect 251646 507922 251702 507978
rect 251274 490294 251330 490350
rect 251398 490294 251454 490350
rect 251522 490294 251578 490350
rect 251646 490294 251702 490350
rect 251274 490170 251330 490226
rect 251398 490170 251454 490226
rect 251522 490170 251578 490226
rect 251646 490170 251702 490226
rect 251274 490046 251330 490102
rect 251398 490046 251454 490102
rect 251522 490046 251578 490102
rect 251646 490046 251702 490102
rect 251274 489922 251330 489978
rect 251398 489922 251454 489978
rect 251522 489922 251578 489978
rect 251646 489922 251702 489978
rect 251274 472294 251330 472350
rect 251398 472294 251454 472350
rect 251522 472294 251578 472350
rect 251646 472294 251702 472350
rect 251274 472170 251330 472226
rect 251398 472170 251454 472226
rect 251522 472170 251578 472226
rect 251646 472170 251702 472226
rect 251274 472046 251330 472102
rect 251398 472046 251454 472102
rect 251522 472046 251578 472102
rect 251646 472046 251702 472102
rect 251274 471922 251330 471978
rect 251398 471922 251454 471978
rect 251522 471922 251578 471978
rect 251646 471922 251702 471978
rect 251274 454294 251330 454350
rect 251398 454294 251454 454350
rect 251522 454294 251578 454350
rect 251646 454294 251702 454350
rect 251274 454170 251330 454226
rect 251398 454170 251454 454226
rect 251522 454170 251578 454226
rect 251646 454170 251702 454226
rect 251274 454046 251330 454102
rect 251398 454046 251454 454102
rect 251522 454046 251578 454102
rect 251646 454046 251702 454102
rect 251274 453922 251330 453978
rect 251398 453922 251454 453978
rect 251522 453922 251578 453978
rect 251646 453922 251702 453978
rect 251274 436294 251330 436350
rect 251398 436294 251454 436350
rect 251522 436294 251578 436350
rect 251646 436294 251702 436350
rect 251274 436170 251330 436226
rect 251398 436170 251454 436226
rect 251522 436170 251578 436226
rect 251646 436170 251702 436226
rect 251274 436046 251330 436102
rect 251398 436046 251454 436102
rect 251522 436046 251578 436102
rect 251646 436046 251702 436102
rect 251274 435922 251330 435978
rect 251398 435922 251454 435978
rect 251522 435922 251578 435978
rect 251646 435922 251702 435978
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 254994 568294 255050 568350
rect 255118 568294 255174 568350
rect 255242 568294 255298 568350
rect 255366 568294 255422 568350
rect 254994 568170 255050 568226
rect 255118 568170 255174 568226
rect 255242 568170 255298 568226
rect 255366 568170 255422 568226
rect 254994 568046 255050 568102
rect 255118 568046 255174 568102
rect 255242 568046 255298 568102
rect 255366 568046 255422 568102
rect 254994 567922 255050 567978
rect 255118 567922 255174 567978
rect 255242 567922 255298 567978
rect 255366 567922 255422 567978
rect 254994 550294 255050 550350
rect 255118 550294 255174 550350
rect 255242 550294 255298 550350
rect 255366 550294 255422 550350
rect 254994 550170 255050 550226
rect 255118 550170 255174 550226
rect 255242 550170 255298 550226
rect 255366 550170 255422 550226
rect 254994 550046 255050 550102
rect 255118 550046 255174 550102
rect 255242 550046 255298 550102
rect 255366 550046 255422 550102
rect 254994 549922 255050 549978
rect 255118 549922 255174 549978
rect 255242 549922 255298 549978
rect 255366 549922 255422 549978
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 281994 562294 282050 562350
rect 282118 562294 282174 562350
rect 282242 562294 282298 562350
rect 282366 562294 282422 562350
rect 281994 562170 282050 562226
rect 282118 562170 282174 562226
rect 282242 562170 282298 562226
rect 282366 562170 282422 562226
rect 281994 562046 282050 562102
rect 282118 562046 282174 562102
rect 282242 562046 282298 562102
rect 282366 562046 282422 562102
rect 281994 561922 282050 561978
rect 282118 561922 282174 561978
rect 282242 561922 282298 561978
rect 282366 561922 282422 561978
rect 268716 546362 268772 546418
rect 254994 532294 255050 532350
rect 255118 532294 255174 532350
rect 255242 532294 255298 532350
rect 255366 532294 255422 532350
rect 254994 532170 255050 532226
rect 255118 532170 255174 532226
rect 255242 532170 255298 532226
rect 255366 532170 255422 532226
rect 254994 532046 255050 532102
rect 255118 532046 255174 532102
rect 255242 532046 255298 532102
rect 255366 532046 255422 532102
rect 254994 531922 255050 531978
rect 255118 531922 255174 531978
rect 255242 531922 255298 531978
rect 255366 531922 255422 531978
rect 254994 514294 255050 514350
rect 255118 514294 255174 514350
rect 255242 514294 255298 514350
rect 255366 514294 255422 514350
rect 254994 514170 255050 514226
rect 255118 514170 255174 514226
rect 255242 514170 255298 514226
rect 255366 514170 255422 514226
rect 254994 514046 255050 514102
rect 255118 514046 255174 514102
rect 255242 514046 255298 514102
rect 255366 514046 255422 514102
rect 254994 513922 255050 513978
rect 255118 513922 255174 513978
rect 255242 513922 255298 513978
rect 255366 513922 255422 513978
rect 254994 496294 255050 496350
rect 255118 496294 255174 496350
rect 255242 496294 255298 496350
rect 255366 496294 255422 496350
rect 254994 496170 255050 496226
rect 255118 496170 255174 496226
rect 255242 496170 255298 496226
rect 255366 496170 255422 496226
rect 254994 496046 255050 496102
rect 255118 496046 255174 496102
rect 255242 496046 255298 496102
rect 255366 496046 255422 496102
rect 254994 495922 255050 495978
rect 255118 495922 255174 495978
rect 255242 495922 255298 495978
rect 255366 495922 255422 495978
rect 254994 478294 255050 478350
rect 255118 478294 255174 478350
rect 255242 478294 255298 478350
rect 255366 478294 255422 478350
rect 254994 478170 255050 478226
rect 255118 478170 255174 478226
rect 255242 478170 255298 478226
rect 255366 478170 255422 478226
rect 254994 478046 255050 478102
rect 255118 478046 255174 478102
rect 255242 478046 255298 478102
rect 255366 478046 255422 478102
rect 254994 477922 255050 477978
rect 255118 477922 255174 477978
rect 255242 477922 255298 477978
rect 255366 477922 255422 477978
rect 254994 460294 255050 460350
rect 255118 460294 255174 460350
rect 255242 460294 255298 460350
rect 255366 460294 255422 460350
rect 254994 460170 255050 460226
rect 255118 460170 255174 460226
rect 255242 460170 255298 460226
rect 255366 460170 255422 460226
rect 254994 460046 255050 460102
rect 255118 460046 255174 460102
rect 255242 460046 255298 460102
rect 255366 460046 255422 460102
rect 254994 459922 255050 459978
rect 255118 459922 255174 459978
rect 255242 459922 255298 459978
rect 255366 459922 255422 459978
rect 254994 442294 255050 442350
rect 255118 442294 255174 442350
rect 255242 442294 255298 442350
rect 255366 442294 255422 442350
rect 254994 442170 255050 442226
rect 255118 442170 255174 442226
rect 255242 442170 255298 442226
rect 255366 442170 255422 442226
rect 254994 442046 255050 442102
rect 255118 442046 255174 442102
rect 255242 442046 255298 442102
rect 255366 442046 255422 442102
rect 254994 441922 255050 441978
rect 255118 441922 255174 441978
rect 255242 441922 255298 441978
rect 255366 441922 255422 441978
rect 267036 546182 267092 546238
rect 281994 544294 282050 544350
rect 282118 544294 282174 544350
rect 282242 544294 282298 544350
rect 282366 544294 282422 544350
rect 281994 544170 282050 544226
rect 282118 544170 282174 544226
rect 282242 544170 282298 544226
rect 282366 544170 282422 544226
rect 281994 544046 282050 544102
rect 282118 544046 282174 544102
rect 282242 544046 282298 544102
rect 282366 544046 282422 544102
rect 281994 543922 282050 543978
rect 282118 543922 282174 543978
rect 282242 543922 282298 543978
rect 282366 543922 282422 543978
rect 281994 526294 282050 526350
rect 282118 526294 282174 526350
rect 282242 526294 282298 526350
rect 282366 526294 282422 526350
rect 281994 526170 282050 526226
rect 282118 526170 282174 526226
rect 282242 526170 282298 526226
rect 282366 526170 282422 526226
rect 281994 526046 282050 526102
rect 282118 526046 282174 526102
rect 282242 526046 282298 526102
rect 282366 526046 282422 526102
rect 281994 525922 282050 525978
rect 282118 525922 282174 525978
rect 282242 525922 282298 525978
rect 282366 525922 282422 525978
rect 281994 508294 282050 508350
rect 282118 508294 282174 508350
rect 282242 508294 282298 508350
rect 282366 508294 282422 508350
rect 281994 508170 282050 508226
rect 282118 508170 282174 508226
rect 282242 508170 282298 508226
rect 282366 508170 282422 508226
rect 281994 508046 282050 508102
rect 282118 508046 282174 508102
rect 282242 508046 282298 508102
rect 282366 508046 282422 508102
rect 281994 507922 282050 507978
rect 282118 507922 282174 507978
rect 282242 507922 282298 507978
rect 282366 507922 282422 507978
rect 281994 490294 282050 490350
rect 282118 490294 282174 490350
rect 282242 490294 282298 490350
rect 282366 490294 282422 490350
rect 281994 490170 282050 490226
rect 282118 490170 282174 490226
rect 282242 490170 282298 490226
rect 282366 490170 282422 490226
rect 281994 490046 282050 490102
rect 282118 490046 282174 490102
rect 282242 490046 282298 490102
rect 282366 490046 282422 490102
rect 281994 489922 282050 489978
rect 282118 489922 282174 489978
rect 282242 489922 282298 489978
rect 282366 489922 282422 489978
rect 281994 472294 282050 472350
rect 282118 472294 282174 472350
rect 282242 472294 282298 472350
rect 282366 472294 282422 472350
rect 281994 472170 282050 472226
rect 282118 472170 282174 472226
rect 282242 472170 282298 472226
rect 282366 472170 282422 472226
rect 281994 472046 282050 472102
rect 282118 472046 282174 472102
rect 282242 472046 282298 472102
rect 282366 472046 282422 472102
rect 281994 471922 282050 471978
rect 282118 471922 282174 471978
rect 282242 471922 282298 471978
rect 282366 471922 282422 471978
rect 281994 454294 282050 454350
rect 282118 454294 282174 454350
rect 282242 454294 282298 454350
rect 282366 454294 282422 454350
rect 281994 454170 282050 454226
rect 282118 454170 282174 454226
rect 282242 454170 282298 454226
rect 282366 454170 282422 454226
rect 281994 454046 282050 454102
rect 282118 454046 282174 454102
rect 282242 454046 282298 454102
rect 282366 454046 282422 454102
rect 281994 453922 282050 453978
rect 282118 453922 282174 453978
rect 282242 453922 282298 453978
rect 282366 453922 282422 453978
rect 281994 436294 282050 436350
rect 282118 436294 282174 436350
rect 282242 436294 282298 436350
rect 282366 436294 282422 436350
rect 281994 436170 282050 436226
rect 282118 436170 282174 436226
rect 282242 436170 282298 436226
rect 282366 436170 282422 436226
rect 281994 436046 282050 436102
rect 282118 436046 282174 436102
rect 282242 436046 282298 436102
rect 282366 436046 282422 436102
rect 281994 435922 282050 435978
rect 282118 435922 282174 435978
rect 282242 435922 282298 435978
rect 282366 435922 282422 435978
rect 276332 432062 276388 432118
rect 110598 424294 110654 424350
rect 110722 424294 110778 424350
rect 110598 424170 110654 424226
rect 110722 424170 110778 424226
rect 110598 424046 110654 424102
rect 110722 424046 110778 424102
rect 110598 423922 110654 423978
rect 110722 423922 110778 423978
rect 141318 424294 141374 424350
rect 141442 424294 141498 424350
rect 141318 424170 141374 424226
rect 141442 424170 141498 424226
rect 141318 424046 141374 424102
rect 141442 424046 141498 424102
rect 141318 423922 141374 423978
rect 141442 423922 141498 423978
rect 172038 424294 172094 424350
rect 172162 424294 172218 424350
rect 172038 424170 172094 424226
rect 172162 424170 172218 424226
rect 172038 424046 172094 424102
rect 172162 424046 172218 424102
rect 172038 423922 172094 423978
rect 172162 423922 172218 423978
rect 202758 424294 202814 424350
rect 202882 424294 202938 424350
rect 202758 424170 202814 424226
rect 202882 424170 202938 424226
rect 202758 424046 202814 424102
rect 202882 424046 202938 424102
rect 202758 423922 202814 423978
rect 202882 423922 202938 423978
rect 233478 424294 233534 424350
rect 233602 424294 233658 424350
rect 233478 424170 233534 424226
rect 233602 424170 233658 424226
rect 233478 424046 233534 424102
rect 233602 424046 233658 424102
rect 233478 423922 233534 423978
rect 233602 423922 233658 423978
rect 95238 418294 95294 418350
rect 95362 418294 95418 418350
rect 95238 418170 95294 418226
rect 95362 418170 95418 418226
rect 95238 418046 95294 418102
rect 95362 418046 95418 418102
rect 95238 417922 95294 417978
rect 95362 417922 95418 417978
rect 125958 418294 126014 418350
rect 126082 418294 126138 418350
rect 125958 418170 126014 418226
rect 126082 418170 126138 418226
rect 125958 418046 126014 418102
rect 126082 418046 126138 418102
rect 125958 417922 126014 417978
rect 126082 417922 126138 417978
rect 156678 418294 156734 418350
rect 156802 418294 156858 418350
rect 156678 418170 156734 418226
rect 156802 418170 156858 418226
rect 156678 418046 156734 418102
rect 156802 418046 156858 418102
rect 156678 417922 156734 417978
rect 156802 417922 156858 417978
rect 187398 418294 187454 418350
rect 187522 418294 187578 418350
rect 187398 418170 187454 418226
rect 187522 418170 187578 418226
rect 187398 418046 187454 418102
rect 187522 418046 187578 418102
rect 187398 417922 187454 417978
rect 187522 417922 187578 417978
rect 218118 418294 218174 418350
rect 218242 418294 218298 418350
rect 218118 418170 218174 418226
rect 218242 418170 218298 418226
rect 218118 418046 218174 418102
rect 218242 418046 218298 418102
rect 218118 417922 218174 417978
rect 218242 417922 218298 417978
rect 248838 418294 248894 418350
rect 248962 418294 249018 418350
rect 248838 418170 248894 418226
rect 248962 418170 249018 418226
rect 248838 418046 248894 418102
rect 248962 418046 249018 418102
rect 248838 417922 248894 417978
rect 248962 417922 249018 417978
rect 83580 409742 83636 409798
rect 110598 406294 110654 406350
rect 110722 406294 110778 406350
rect 110598 406170 110654 406226
rect 110722 406170 110778 406226
rect 110598 406046 110654 406102
rect 110722 406046 110778 406102
rect 110598 405922 110654 405978
rect 110722 405922 110778 405978
rect 141318 406294 141374 406350
rect 141442 406294 141498 406350
rect 141318 406170 141374 406226
rect 141442 406170 141498 406226
rect 141318 406046 141374 406102
rect 141442 406046 141498 406102
rect 141318 405922 141374 405978
rect 141442 405922 141498 405978
rect 172038 406294 172094 406350
rect 172162 406294 172218 406350
rect 172038 406170 172094 406226
rect 172162 406170 172218 406226
rect 172038 406046 172094 406102
rect 172162 406046 172218 406102
rect 172038 405922 172094 405978
rect 172162 405922 172218 405978
rect 202758 406294 202814 406350
rect 202882 406294 202938 406350
rect 202758 406170 202814 406226
rect 202882 406170 202938 406226
rect 202758 406046 202814 406102
rect 202882 406046 202938 406102
rect 202758 405922 202814 405978
rect 202882 405922 202938 405978
rect 233478 406294 233534 406350
rect 233602 406294 233658 406350
rect 233478 406170 233534 406226
rect 233602 406170 233658 406226
rect 233478 406046 233534 406102
rect 233602 406046 233658 406102
rect 233478 405922 233534 405978
rect 233602 405922 233658 405978
rect 260316 403082 260372 403138
rect 264198 424294 264254 424350
rect 264322 424294 264378 424350
rect 264198 424170 264254 424226
rect 264322 424170 264378 424226
rect 264198 424046 264254 424102
rect 264322 424046 264378 424102
rect 264198 423922 264254 423978
rect 264322 423922 264378 423978
rect 264198 406294 264254 406350
rect 264322 406294 264378 406350
rect 264198 406170 264254 406226
rect 264322 406170 264378 406226
rect 264198 406046 264254 406102
rect 264322 406046 264378 406102
rect 264198 405922 264254 405978
rect 264322 405922 264378 405978
rect 263676 402902 263732 402958
rect 95238 400294 95294 400350
rect 95362 400294 95418 400350
rect 95238 400170 95294 400226
rect 95362 400170 95418 400226
rect 95238 400046 95294 400102
rect 95362 400046 95418 400102
rect 95238 399922 95294 399978
rect 95362 399922 95418 399978
rect 125958 400294 126014 400350
rect 126082 400294 126138 400350
rect 125958 400170 126014 400226
rect 126082 400170 126138 400226
rect 125958 400046 126014 400102
rect 126082 400046 126138 400102
rect 125958 399922 126014 399978
rect 126082 399922 126138 399978
rect 156678 400294 156734 400350
rect 156802 400294 156858 400350
rect 156678 400170 156734 400226
rect 156802 400170 156858 400226
rect 156678 400046 156734 400102
rect 156802 400046 156858 400102
rect 156678 399922 156734 399978
rect 156802 399922 156858 399978
rect 187398 400294 187454 400350
rect 187522 400294 187578 400350
rect 187398 400170 187454 400226
rect 187522 400170 187578 400226
rect 187398 400046 187454 400102
rect 187522 400046 187578 400102
rect 187398 399922 187454 399978
rect 187522 399922 187578 399978
rect 218118 400294 218174 400350
rect 218242 400294 218298 400350
rect 218118 400170 218174 400226
rect 218242 400170 218298 400226
rect 218118 400046 218174 400102
rect 218242 400046 218298 400102
rect 218118 399922 218174 399978
rect 218242 399922 218298 399978
rect 248838 400294 248894 400350
rect 248962 400294 249018 400350
rect 248838 400170 248894 400226
rect 248962 400170 249018 400226
rect 248838 400046 248894 400102
rect 248962 400046 249018 400102
rect 248838 399922 248894 399978
rect 248962 399922 249018 399978
rect 110598 388294 110654 388350
rect 110722 388294 110778 388350
rect 110598 388170 110654 388226
rect 110722 388170 110778 388226
rect 110598 388046 110654 388102
rect 110722 388046 110778 388102
rect 110598 387922 110654 387978
rect 110722 387922 110778 387978
rect 141318 388294 141374 388350
rect 141442 388294 141498 388350
rect 141318 388170 141374 388226
rect 141442 388170 141498 388226
rect 141318 388046 141374 388102
rect 141442 388046 141498 388102
rect 141318 387922 141374 387978
rect 141442 387922 141498 387978
rect 172038 388294 172094 388350
rect 172162 388294 172218 388350
rect 172038 388170 172094 388226
rect 172162 388170 172218 388226
rect 172038 388046 172094 388102
rect 172162 388046 172218 388102
rect 172038 387922 172094 387978
rect 172162 387922 172218 387978
rect 202758 388294 202814 388350
rect 202882 388294 202938 388350
rect 202758 388170 202814 388226
rect 202882 388170 202938 388226
rect 202758 388046 202814 388102
rect 202882 388046 202938 388102
rect 202758 387922 202814 387978
rect 202882 387922 202938 387978
rect 233478 388294 233534 388350
rect 233602 388294 233658 388350
rect 233478 388170 233534 388226
rect 233602 388170 233658 388226
rect 233478 388046 233534 388102
rect 233602 388046 233658 388102
rect 233478 387922 233534 387978
rect 233602 387922 233658 387978
rect 264198 388294 264254 388350
rect 264322 388294 264378 388350
rect 264198 388170 264254 388226
rect 264322 388170 264378 388226
rect 264198 388046 264254 388102
rect 264322 388046 264378 388102
rect 264198 387922 264254 387978
rect 264322 387922 264378 387978
rect 84812 383102 84868 383158
rect 83468 347642 83524 347698
rect 83580 368162 83636 368218
rect 83804 367982 83860 368038
rect 83580 295262 83636 295318
rect 83692 366362 83748 366418
rect 95238 382294 95294 382350
rect 95362 382294 95418 382350
rect 95238 382170 95294 382226
rect 95362 382170 95418 382226
rect 95238 382046 95294 382102
rect 95362 382046 95418 382102
rect 95238 381922 95294 381978
rect 95362 381922 95418 381978
rect 125958 382294 126014 382350
rect 126082 382294 126138 382350
rect 125958 382170 126014 382226
rect 126082 382170 126138 382226
rect 125958 382046 126014 382102
rect 126082 382046 126138 382102
rect 125958 381922 126014 381978
rect 126082 381922 126138 381978
rect 156678 382294 156734 382350
rect 156802 382294 156858 382350
rect 156678 382170 156734 382226
rect 156802 382170 156858 382226
rect 156678 382046 156734 382102
rect 156802 382046 156858 382102
rect 156678 381922 156734 381978
rect 156802 381922 156858 381978
rect 187398 382294 187454 382350
rect 187522 382294 187578 382350
rect 187398 382170 187454 382226
rect 187522 382170 187578 382226
rect 187398 382046 187454 382102
rect 187522 382046 187578 382102
rect 187398 381922 187454 381978
rect 187522 381922 187578 381978
rect 218118 382294 218174 382350
rect 218242 382294 218298 382350
rect 218118 382170 218174 382226
rect 218242 382170 218298 382226
rect 218118 382046 218174 382102
rect 218242 382046 218298 382102
rect 218118 381922 218174 381978
rect 218242 381922 218298 381978
rect 248838 382294 248894 382350
rect 248962 382294 249018 382350
rect 248838 382170 248894 382226
rect 248962 382170 249018 382226
rect 248838 382046 248894 382102
rect 248962 382046 249018 382102
rect 273532 388862 273588 388918
rect 248838 381922 248894 381978
rect 248962 381922 249018 381978
rect 276444 387602 276500 387658
rect 273756 371402 273812 371458
rect 110598 370294 110654 370350
rect 110722 370294 110778 370350
rect 110598 370170 110654 370226
rect 110722 370170 110778 370226
rect 110598 370046 110654 370102
rect 110722 370046 110778 370102
rect 110598 369922 110654 369978
rect 110722 369922 110778 369978
rect 141318 370294 141374 370350
rect 141442 370294 141498 370350
rect 141318 370170 141374 370226
rect 141442 370170 141498 370226
rect 141318 370046 141374 370102
rect 141442 370046 141498 370102
rect 141318 369922 141374 369978
rect 141442 369922 141498 369978
rect 172038 370294 172094 370350
rect 172162 370294 172218 370350
rect 172038 370170 172094 370226
rect 172162 370170 172218 370226
rect 172038 370046 172094 370102
rect 172162 370046 172218 370102
rect 172038 369922 172094 369978
rect 172162 369922 172218 369978
rect 202758 370294 202814 370350
rect 202882 370294 202938 370350
rect 202758 370170 202814 370226
rect 202882 370170 202938 370226
rect 202758 370046 202814 370102
rect 202882 370046 202938 370102
rect 202758 369922 202814 369978
rect 202882 369922 202938 369978
rect 233478 370294 233534 370350
rect 233602 370294 233658 370350
rect 233478 370170 233534 370226
rect 233602 370170 233658 370226
rect 233478 370046 233534 370102
rect 233602 370046 233658 370102
rect 233478 369922 233534 369978
rect 233602 369922 233658 369978
rect 264198 370294 264254 370350
rect 264322 370294 264378 370350
rect 264198 370170 264254 370226
rect 264322 370170 264378 370226
rect 264198 370046 264254 370102
rect 264322 370046 264378 370102
rect 264198 369922 264254 369978
rect 264322 369922 264378 369978
rect 273756 367982 273812 368038
rect 273756 366362 273812 366418
rect 273756 364742 273812 364798
rect 273756 364588 273812 364618
rect 273756 364562 273812 364588
rect 95238 364294 95294 364350
rect 95362 364294 95418 364350
rect 95238 364170 95294 364226
rect 95362 364170 95418 364226
rect 95238 364046 95294 364102
rect 95362 364046 95418 364102
rect 95238 363922 95294 363978
rect 95362 363922 95418 363978
rect 125958 364294 126014 364350
rect 126082 364294 126138 364350
rect 125958 364170 126014 364226
rect 126082 364170 126138 364226
rect 125958 364046 126014 364102
rect 126082 364046 126138 364102
rect 125958 363922 126014 363978
rect 126082 363922 126138 363978
rect 156678 364294 156734 364350
rect 156802 364294 156858 364350
rect 156678 364170 156734 364226
rect 156802 364170 156858 364226
rect 156678 364046 156734 364102
rect 156802 364046 156858 364102
rect 156678 363922 156734 363978
rect 156802 363922 156858 363978
rect 187398 364294 187454 364350
rect 187522 364294 187578 364350
rect 187398 364170 187454 364226
rect 187522 364170 187578 364226
rect 187398 364046 187454 364102
rect 187522 364046 187578 364102
rect 187398 363922 187454 363978
rect 187522 363922 187578 363978
rect 218118 364294 218174 364350
rect 218242 364294 218298 364350
rect 218118 364170 218174 364226
rect 218242 364170 218298 364226
rect 218118 364046 218174 364102
rect 218242 364046 218298 364102
rect 218118 363922 218174 363978
rect 218242 363922 218298 363978
rect 248838 364294 248894 364350
rect 248962 364294 249018 364350
rect 248838 364170 248894 364226
rect 248962 364170 249018 364226
rect 248838 364046 248894 364102
rect 248962 364046 249018 364102
rect 248838 363922 248894 363978
rect 248962 363922 249018 363978
rect 110598 352294 110654 352350
rect 110722 352294 110778 352350
rect 110598 352170 110654 352226
rect 110722 352170 110778 352226
rect 110598 352046 110654 352102
rect 110722 352046 110778 352102
rect 110598 351922 110654 351978
rect 110722 351922 110778 351978
rect 141318 352294 141374 352350
rect 141442 352294 141498 352350
rect 141318 352170 141374 352226
rect 141442 352170 141498 352226
rect 141318 352046 141374 352102
rect 141442 352046 141498 352102
rect 141318 351922 141374 351978
rect 141442 351922 141498 351978
rect 172038 352294 172094 352350
rect 172162 352294 172218 352350
rect 172038 352170 172094 352226
rect 172162 352170 172218 352226
rect 172038 352046 172094 352102
rect 172162 352046 172218 352102
rect 172038 351922 172094 351978
rect 172162 351922 172218 351978
rect 202758 352294 202814 352350
rect 202882 352294 202938 352350
rect 202758 352170 202814 352226
rect 202882 352170 202938 352226
rect 202758 352046 202814 352102
rect 202882 352046 202938 352102
rect 202758 351922 202814 351978
rect 202882 351922 202938 351978
rect 233478 352294 233534 352350
rect 233602 352294 233658 352350
rect 233478 352170 233534 352226
rect 233602 352170 233658 352226
rect 233478 352046 233534 352102
rect 233602 352046 233658 352102
rect 233478 351922 233534 351978
rect 233602 351922 233658 351978
rect 264198 352294 264254 352350
rect 264322 352294 264378 352350
rect 264198 352170 264254 352226
rect 264322 352170 264378 352226
rect 264198 352046 264254 352102
rect 264322 352046 264378 352102
rect 264198 351922 264254 351978
rect 264322 351922 264378 351978
rect 95238 346294 95294 346350
rect 95362 346294 95418 346350
rect 95238 346170 95294 346226
rect 95362 346170 95418 346226
rect 95238 346046 95294 346102
rect 95362 346046 95418 346102
rect 95238 345922 95294 345978
rect 95362 345922 95418 345978
rect 125958 346294 126014 346350
rect 126082 346294 126138 346350
rect 125958 346170 126014 346226
rect 126082 346170 126138 346226
rect 125958 346046 126014 346102
rect 126082 346046 126138 346102
rect 125958 345922 126014 345978
rect 126082 345922 126138 345978
rect 156678 346294 156734 346350
rect 156802 346294 156858 346350
rect 156678 346170 156734 346226
rect 156802 346170 156858 346226
rect 156678 346046 156734 346102
rect 156802 346046 156858 346102
rect 156678 345922 156734 345978
rect 156802 345922 156858 345978
rect 187398 346294 187454 346350
rect 187522 346294 187578 346350
rect 187398 346170 187454 346226
rect 187522 346170 187578 346226
rect 187398 346046 187454 346102
rect 187522 346046 187578 346102
rect 187398 345922 187454 345978
rect 187522 345922 187578 345978
rect 218118 346294 218174 346350
rect 218242 346294 218298 346350
rect 218118 346170 218174 346226
rect 218242 346170 218298 346226
rect 218118 346046 218174 346102
rect 218242 346046 218298 346102
rect 218118 345922 218174 345978
rect 218242 345922 218298 345978
rect 248838 346294 248894 346350
rect 248962 346294 249018 346350
rect 248838 346170 248894 346226
rect 248962 346170 249018 346226
rect 248838 346046 248894 346102
rect 248962 346046 249018 346102
rect 248838 345922 248894 345978
rect 248962 345922 249018 345978
rect 110598 334294 110654 334350
rect 110722 334294 110778 334350
rect 110598 334170 110654 334226
rect 110722 334170 110778 334226
rect 110598 334046 110654 334102
rect 110722 334046 110778 334102
rect 110598 333922 110654 333978
rect 110722 333922 110778 333978
rect 141318 334294 141374 334350
rect 141442 334294 141498 334350
rect 141318 334170 141374 334226
rect 141442 334170 141498 334226
rect 141318 334046 141374 334102
rect 141442 334046 141498 334102
rect 141318 333922 141374 333978
rect 141442 333922 141498 333978
rect 172038 334294 172094 334350
rect 172162 334294 172218 334350
rect 172038 334170 172094 334226
rect 172162 334170 172218 334226
rect 172038 334046 172094 334102
rect 172162 334046 172218 334102
rect 172038 333922 172094 333978
rect 172162 333922 172218 333978
rect 202758 334294 202814 334350
rect 202882 334294 202938 334350
rect 202758 334170 202814 334226
rect 202882 334170 202938 334226
rect 202758 334046 202814 334102
rect 202882 334046 202938 334102
rect 202758 333922 202814 333978
rect 202882 333922 202938 333978
rect 233478 334294 233534 334350
rect 233602 334294 233658 334350
rect 233478 334170 233534 334226
rect 233602 334170 233658 334226
rect 233478 334046 233534 334102
rect 233602 334046 233658 334102
rect 233478 333922 233534 333978
rect 233602 333922 233658 333978
rect 264198 334294 264254 334350
rect 264322 334294 264378 334350
rect 264198 334170 264254 334226
rect 264322 334170 264378 334226
rect 264198 334046 264254 334102
rect 264322 334046 264378 334102
rect 264198 333922 264254 333978
rect 264322 333922 264378 333978
rect 84812 300122 84868 300178
rect 84924 329282 84980 329338
rect 83804 298862 83860 298918
rect 95238 328294 95294 328350
rect 95362 328294 95418 328350
rect 95238 328170 95294 328226
rect 95362 328170 95418 328226
rect 95238 328046 95294 328102
rect 95362 328046 95418 328102
rect 95238 327922 95294 327978
rect 95362 327922 95418 327978
rect 125958 328294 126014 328350
rect 126082 328294 126138 328350
rect 125958 328170 126014 328226
rect 126082 328170 126138 328226
rect 125958 328046 126014 328102
rect 126082 328046 126138 328102
rect 125958 327922 126014 327978
rect 126082 327922 126138 327978
rect 156678 328294 156734 328350
rect 156802 328294 156858 328350
rect 156678 328170 156734 328226
rect 156802 328170 156858 328226
rect 156678 328046 156734 328102
rect 156802 328046 156858 328102
rect 156678 327922 156734 327978
rect 156802 327922 156858 327978
rect 187398 328294 187454 328350
rect 187522 328294 187578 328350
rect 187398 328170 187454 328226
rect 187522 328170 187578 328226
rect 187398 328046 187454 328102
rect 187522 328046 187578 328102
rect 187398 327922 187454 327978
rect 187522 327922 187578 327978
rect 218118 328294 218174 328350
rect 218242 328294 218298 328350
rect 218118 328170 218174 328226
rect 218242 328170 218298 328226
rect 218118 328046 218174 328102
rect 218242 328046 218298 328102
rect 218118 327922 218174 327978
rect 218242 327922 218298 327978
rect 248838 328294 248894 328350
rect 248962 328294 249018 328350
rect 248838 328170 248894 328226
rect 248962 328170 249018 328226
rect 248838 328046 248894 328102
rect 248962 328046 249018 328102
rect 248838 327922 248894 327978
rect 248962 327922 249018 327978
rect 273756 361322 273812 361378
rect 273756 358622 273812 358678
rect 273756 356282 273812 356338
rect 273756 354482 273812 354538
rect 273756 353582 273812 353638
rect 273308 350162 273364 350218
rect 273084 343502 273140 343558
rect 273756 349442 273812 349498
rect 273756 343682 273812 343738
rect 273644 341882 273700 341938
rect 272972 319922 273028 319978
rect 110598 316294 110654 316350
rect 110722 316294 110778 316350
rect 110598 316170 110654 316226
rect 110722 316170 110778 316226
rect 110598 316046 110654 316102
rect 110722 316046 110778 316102
rect 110598 315922 110654 315978
rect 110722 315922 110778 315978
rect 141318 316294 141374 316350
rect 141442 316294 141498 316350
rect 141318 316170 141374 316226
rect 141442 316170 141498 316226
rect 141318 316046 141374 316102
rect 141442 316046 141498 316102
rect 141318 315922 141374 315978
rect 141442 315922 141498 315978
rect 172038 316294 172094 316350
rect 172162 316294 172218 316350
rect 172038 316170 172094 316226
rect 172162 316170 172218 316226
rect 172038 316046 172094 316102
rect 172162 316046 172218 316102
rect 172038 315922 172094 315978
rect 172162 315922 172218 315978
rect 202758 316294 202814 316350
rect 202882 316294 202938 316350
rect 202758 316170 202814 316226
rect 202882 316170 202938 316226
rect 202758 316046 202814 316102
rect 202882 316046 202938 316102
rect 202758 315922 202814 315978
rect 202882 315922 202938 315978
rect 233478 316294 233534 316350
rect 233602 316294 233658 316350
rect 233478 316170 233534 316226
rect 233602 316170 233658 316226
rect 233478 316046 233534 316102
rect 233602 316046 233658 316102
rect 233478 315922 233534 315978
rect 233602 315922 233658 315978
rect 264198 316294 264254 316350
rect 264322 316294 264378 316350
rect 264198 316170 264254 316226
rect 264322 316170 264378 316226
rect 264198 316046 264254 316102
rect 264322 316046 264378 316102
rect 264198 315922 264254 315978
rect 264322 315922 264378 315978
rect 278124 335942 278180 335998
rect 278236 376442 278292 376498
rect 278012 333602 278068 333658
rect 273756 330002 273812 330058
rect 273308 324962 273364 325018
rect 273196 323342 273252 323398
rect 273084 311642 273140 311698
rect 274652 317582 274708 317638
rect 95238 310294 95294 310350
rect 95362 310294 95418 310350
rect 95238 310170 95294 310226
rect 95362 310170 95418 310226
rect 95238 310046 95294 310102
rect 95362 310046 95418 310102
rect 95238 309922 95294 309978
rect 95362 309922 95418 309978
rect 125958 310294 126014 310350
rect 126082 310294 126138 310350
rect 125958 310170 126014 310226
rect 126082 310170 126138 310226
rect 125958 310046 126014 310102
rect 126082 310046 126138 310102
rect 125958 309922 126014 309978
rect 126082 309922 126138 309978
rect 156678 310294 156734 310350
rect 156802 310294 156858 310350
rect 156678 310170 156734 310226
rect 156802 310170 156858 310226
rect 156678 310046 156734 310102
rect 156802 310046 156858 310102
rect 156678 309922 156734 309978
rect 156802 309922 156858 309978
rect 187398 310294 187454 310350
rect 187522 310294 187578 310350
rect 187398 310170 187454 310226
rect 187522 310170 187578 310226
rect 187398 310046 187454 310102
rect 187522 310046 187578 310102
rect 187398 309922 187454 309978
rect 187522 309922 187578 309978
rect 218118 310294 218174 310350
rect 218242 310294 218298 310350
rect 218118 310170 218174 310226
rect 218242 310170 218298 310226
rect 218118 310046 218174 310102
rect 218242 310046 218298 310102
rect 218118 309922 218174 309978
rect 218242 309922 218298 309978
rect 248838 310294 248894 310350
rect 248962 310294 249018 310350
rect 248838 310170 248894 310226
rect 248962 310170 249018 310226
rect 248838 310046 248894 310102
rect 248962 310046 249018 310102
rect 248838 309922 248894 309978
rect 248962 309922 249018 309978
rect 84924 297242 84980 297298
rect 83692 295082 83748 295138
rect 97674 292294 97730 292350
rect 97798 292294 97854 292350
rect 97922 292294 97978 292350
rect 98046 292294 98102 292350
rect 97674 292170 97730 292226
rect 97798 292170 97854 292226
rect 97922 292170 97978 292226
rect 98046 292170 98102 292226
rect 97674 292046 97730 292102
rect 97798 292046 97854 292102
rect 97922 292046 97978 292102
rect 98046 292046 98102 292102
rect 97674 291922 97730 291978
rect 97798 291922 97854 291978
rect 97922 291922 97978 291978
rect 98046 291922 98102 291978
rect 97674 274294 97730 274350
rect 97798 274294 97854 274350
rect 97922 274294 97978 274350
rect 98046 274294 98102 274350
rect 97674 274170 97730 274226
rect 97798 274170 97854 274226
rect 97922 274170 97978 274226
rect 98046 274170 98102 274226
rect 97674 274046 97730 274102
rect 97798 274046 97854 274102
rect 97922 274046 97978 274102
rect 98046 274046 98102 274102
rect 97674 273922 97730 273978
rect 97798 273922 97854 273978
rect 97922 273922 97978 273978
rect 98046 273922 98102 273978
rect 84924 142082 84980 142138
rect 97674 256294 97730 256350
rect 97798 256294 97854 256350
rect 97922 256294 97978 256350
rect 98046 256294 98102 256350
rect 97674 256170 97730 256226
rect 97798 256170 97854 256226
rect 97922 256170 97978 256226
rect 98046 256170 98102 256226
rect 97674 256046 97730 256102
rect 97798 256046 97854 256102
rect 97922 256046 97978 256102
rect 98046 256046 98102 256102
rect 97674 255922 97730 255978
rect 97798 255922 97854 255978
rect 97922 255922 97978 255978
rect 98046 255922 98102 255978
rect 97674 238294 97730 238350
rect 97798 238294 97854 238350
rect 97922 238294 97978 238350
rect 98046 238294 98102 238350
rect 97674 238170 97730 238226
rect 97798 238170 97854 238226
rect 97922 238170 97978 238226
rect 98046 238170 98102 238226
rect 97674 238046 97730 238102
rect 97798 238046 97854 238102
rect 97922 238046 97978 238102
rect 98046 238046 98102 238102
rect 97674 237922 97730 237978
rect 97798 237922 97854 237978
rect 97922 237922 97978 237978
rect 98046 237922 98102 237978
rect 97674 220294 97730 220350
rect 97798 220294 97854 220350
rect 97922 220294 97978 220350
rect 98046 220294 98102 220350
rect 97674 220170 97730 220226
rect 97798 220170 97854 220226
rect 97922 220170 97978 220226
rect 98046 220170 98102 220226
rect 97674 220046 97730 220102
rect 97798 220046 97854 220102
rect 97922 220046 97978 220102
rect 98046 220046 98102 220102
rect 97674 219922 97730 219978
rect 97798 219922 97854 219978
rect 97922 219922 97978 219978
rect 98046 219922 98102 219978
rect 95238 202294 95294 202350
rect 95362 202294 95418 202350
rect 95238 202170 95294 202226
rect 95362 202170 95418 202226
rect 95238 202046 95294 202102
rect 95362 202046 95418 202102
rect 95238 201922 95294 201978
rect 95362 201922 95418 201978
rect 97674 202294 97730 202350
rect 97798 202294 97854 202350
rect 97922 202294 97978 202350
rect 98046 202294 98102 202350
rect 97674 202170 97730 202226
rect 97798 202170 97854 202226
rect 97922 202170 97978 202226
rect 98046 202170 98102 202226
rect 97674 202046 97730 202102
rect 97798 202046 97854 202102
rect 97922 202046 97978 202102
rect 98046 202046 98102 202102
rect 97674 201922 97730 201978
rect 97798 201922 97854 201978
rect 97922 201922 97978 201978
rect 98046 201922 98102 201978
rect 95238 184294 95294 184350
rect 95362 184294 95418 184350
rect 95238 184170 95294 184226
rect 95362 184170 95418 184226
rect 95238 184046 95294 184102
rect 95362 184046 95418 184102
rect 95238 183922 95294 183978
rect 95362 183922 95418 183978
rect 97674 184294 97730 184350
rect 97798 184294 97854 184350
rect 97922 184294 97978 184350
rect 98046 184294 98102 184350
rect 97674 184170 97730 184226
rect 97798 184170 97854 184226
rect 97922 184170 97978 184226
rect 98046 184170 98102 184226
rect 97674 184046 97730 184102
rect 97798 184046 97854 184102
rect 97922 184046 97978 184102
rect 98046 184046 98102 184102
rect 97674 183922 97730 183978
rect 97798 183922 97854 183978
rect 97922 183922 97978 183978
rect 98046 183922 98102 183978
rect 95238 166294 95294 166350
rect 95362 166294 95418 166350
rect 95238 166170 95294 166226
rect 95362 166170 95418 166226
rect 95238 166046 95294 166102
rect 95362 166046 95418 166102
rect 95238 165922 95294 165978
rect 95362 165922 95418 165978
rect 97674 166294 97730 166350
rect 97798 166294 97854 166350
rect 97922 166294 97978 166350
rect 98046 166294 98102 166350
rect 97674 166170 97730 166226
rect 97798 166170 97854 166226
rect 97922 166170 97978 166226
rect 98046 166170 98102 166226
rect 97674 166046 97730 166102
rect 97798 166046 97854 166102
rect 97922 166046 97978 166102
rect 98046 166046 98102 166102
rect 97674 165922 97730 165978
rect 97798 165922 97854 165978
rect 97922 165922 97978 165978
rect 98046 165922 98102 165978
rect 97674 148294 97730 148350
rect 97798 148294 97854 148350
rect 97922 148294 97978 148350
rect 98046 148294 98102 148350
rect 97674 148170 97730 148226
rect 97798 148170 97854 148226
rect 97922 148170 97978 148226
rect 98046 148170 98102 148226
rect 97674 148046 97730 148102
rect 97798 148046 97854 148102
rect 97922 148046 97978 148102
rect 98046 148046 98102 148102
rect 97674 147922 97730 147978
rect 97798 147922 97854 147978
rect 97922 147922 97978 147978
rect 98046 147922 98102 147978
rect 97674 130294 97730 130350
rect 97798 130294 97854 130350
rect 97922 130294 97978 130350
rect 98046 130294 98102 130350
rect 97674 130170 97730 130226
rect 97798 130170 97854 130226
rect 97922 130170 97978 130226
rect 98046 130170 98102 130226
rect 97674 130046 97730 130102
rect 97798 130046 97854 130102
rect 97922 130046 97978 130102
rect 98046 130046 98102 130102
rect 97674 129922 97730 129978
rect 97798 129922 97854 129978
rect 97922 129922 97978 129978
rect 98046 129922 98102 129978
rect 97674 112294 97730 112350
rect 97798 112294 97854 112350
rect 97922 112294 97978 112350
rect 98046 112294 98102 112350
rect 97674 112170 97730 112226
rect 97798 112170 97854 112226
rect 97922 112170 97978 112226
rect 98046 112170 98102 112226
rect 97674 112046 97730 112102
rect 97798 112046 97854 112102
rect 97922 112046 97978 112102
rect 98046 112046 98102 112102
rect 97674 111922 97730 111978
rect 97798 111922 97854 111978
rect 97922 111922 97978 111978
rect 98046 111922 98102 111978
rect 97674 94294 97730 94350
rect 97798 94294 97854 94350
rect 97922 94294 97978 94350
rect 98046 94294 98102 94350
rect 97674 94170 97730 94226
rect 97798 94170 97854 94226
rect 97922 94170 97978 94226
rect 98046 94170 98102 94226
rect 97674 94046 97730 94102
rect 97798 94046 97854 94102
rect 97922 94046 97978 94102
rect 98046 94046 98102 94102
rect 97674 93922 97730 93978
rect 97798 93922 97854 93978
rect 97922 93922 97978 93978
rect 98046 93922 98102 93978
rect 97674 76294 97730 76350
rect 97798 76294 97854 76350
rect 97922 76294 97978 76350
rect 98046 76294 98102 76350
rect 97674 76170 97730 76226
rect 97798 76170 97854 76226
rect 97922 76170 97978 76226
rect 98046 76170 98102 76226
rect 97674 76046 97730 76102
rect 97798 76046 97854 76102
rect 97922 76046 97978 76102
rect 98046 76046 98102 76102
rect 97674 75922 97730 75978
rect 97798 75922 97854 75978
rect 97922 75922 97978 75978
rect 98046 75922 98102 75978
rect 97674 58294 97730 58350
rect 97798 58294 97854 58350
rect 97922 58294 97978 58350
rect 98046 58294 98102 58350
rect 97674 58170 97730 58226
rect 97798 58170 97854 58226
rect 97922 58170 97978 58226
rect 98046 58170 98102 58226
rect 97674 58046 97730 58102
rect 97798 58046 97854 58102
rect 97922 58046 97978 58102
rect 98046 58046 98102 58102
rect 97674 57922 97730 57978
rect 97798 57922 97854 57978
rect 97922 57922 97978 57978
rect 98046 57922 98102 57978
rect 97674 40294 97730 40350
rect 97798 40294 97854 40350
rect 97922 40294 97978 40350
rect 98046 40294 98102 40350
rect 97674 40170 97730 40226
rect 97798 40170 97854 40226
rect 97922 40170 97978 40226
rect 98046 40170 98102 40226
rect 97674 40046 97730 40102
rect 97798 40046 97854 40102
rect 97922 40046 97978 40102
rect 98046 40046 98102 40102
rect 97674 39922 97730 39978
rect 97798 39922 97854 39978
rect 97922 39922 97978 39978
rect 98046 39922 98102 39978
rect 97674 22294 97730 22350
rect 97798 22294 97854 22350
rect 97922 22294 97978 22350
rect 98046 22294 98102 22350
rect 97674 22170 97730 22226
rect 97798 22170 97854 22226
rect 97922 22170 97978 22226
rect 98046 22170 98102 22226
rect 97674 22046 97730 22102
rect 97798 22046 97854 22102
rect 97922 22046 97978 22102
rect 98046 22046 98102 22102
rect 97674 21922 97730 21978
rect 97798 21922 97854 21978
rect 97922 21922 97978 21978
rect 98046 21922 98102 21978
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 101394 298294 101450 298350
rect 101518 298294 101574 298350
rect 101642 298294 101698 298350
rect 101766 298294 101822 298350
rect 101394 298170 101450 298226
rect 101518 298170 101574 298226
rect 101642 298170 101698 298226
rect 101766 298170 101822 298226
rect 101394 298046 101450 298102
rect 101518 298046 101574 298102
rect 101642 298046 101698 298102
rect 101766 298046 101822 298102
rect 101394 297922 101450 297978
rect 101518 297922 101574 297978
rect 101642 297922 101698 297978
rect 101766 297922 101822 297978
rect 110598 298294 110654 298350
rect 110722 298294 110778 298350
rect 110598 298170 110654 298226
rect 110722 298170 110778 298226
rect 110598 298046 110654 298102
rect 110722 298046 110778 298102
rect 110598 297922 110654 297978
rect 110722 297922 110778 297978
rect 128394 292294 128450 292350
rect 128518 292294 128574 292350
rect 128642 292294 128698 292350
rect 128766 292294 128822 292350
rect 128394 292170 128450 292226
rect 128518 292170 128574 292226
rect 128642 292170 128698 292226
rect 128766 292170 128822 292226
rect 128394 292046 128450 292102
rect 128518 292046 128574 292102
rect 128642 292046 128698 292102
rect 128766 292046 128822 292102
rect 128394 291922 128450 291978
rect 128518 291922 128574 291978
rect 128642 291922 128698 291978
rect 128766 291922 128822 291978
rect 101394 280294 101450 280350
rect 101518 280294 101574 280350
rect 101642 280294 101698 280350
rect 101766 280294 101822 280350
rect 101394 280170 101450 280226
rect 101518 280170 101574 280226
rect 101642 280170 101698 280226
rect 101766 280170 101822 280226
rect 101394 280046 101450 280102
rect 101518 280046 101574 280102
rect 101642 280046 101698 280102
rect 101766 280046 101822 280102
rect 101394 279922 101450 279978
rect 101518 279922 101574 279978
rect 101642 279922 101698 279978
rect 101766 279922 101822 279978
rect 101394 262294 101450 262350
rect 101518 262294 101574 262350
rect 101642 262294 101698 262350
rect 101766 262294 101822 262350
rect 101394 262170 101450 262226
rect 101518 262170 101574 262226
rect 101642 262170 101698 262226
rect 101766 262170 101822 262226
rect 101394 262046 101450 262102
rect 101518 262046 101574 262102
rect 101642 262046 101698 262102
rect 101766 262046 101822 262102
rect 101394 261922 101450 261978
rect 101518 261922 101574 261978
rect 101642 261922 101698 261978
rect 101766 261922 101822 261978
rect 101394 244294 101450 244350
rect 101518 244294 101574 244350
rect 101642 244294 101698 244350
rect 101766 244294 101822 244350
rect 101394 244170 101450 244226
rect 101518 244170 101574 244226
rect 101642 244170 101698 244226
rect 101766 244170 101822 244226
rect 101394 244046 101450 244102
rect 101518 244046 101574 244102
rect 101642 244046 101698 244102
rect 101766 244046 101822 244102
rect 101394 243922 101450 243978
rect 101518 243922 101574 243978
rect 101642 243922 101698 243978
rect 101766 243922 101822 243978
rect 101394 226294 101450 226350
rect 101518 226294 101574 226350
rect 101642 226294 101698 226350
rect 101766 226294 101822 226350
rect 101394 226170 101450 226226
rect 101518 226170 101574 226226
rect 101642 226170 101698 226226
rect 101766 226170 101822 226226
rect 101394 226046 101450 226102
rect 101518 226046 101574 226102
rect 101642 226046 101698 226102
rect 101766 226046 101822 226102
rect 101394 225922 101450 225978
rect 101518 225922 101574 225978
rect 101642 225922 101698 225978
rect 101766 225922 101822 225978
rect 101394 208294 101450 208350
rect 101518 208294 101574 208350
rect 101642 208294 101698 208350
rect 101766 208294 101822 208350
rect 101394 208170 101450 208226
rect 101518 208170 101574 208226
rect 101642 208170 101698 208226
rect 101766 208170 101822 208226
rect 101394 208046 101450 208102
rect 101518 208046 101574 208102
rect 101642 208046 101698 208102
rect 101766 208046 101822 208102
rect 101394 207922 101450 207978
rect 101518 207922 101574 207978
rect 101642 207922 101698 207978
rect 101766 207922 101822 207978
rect 101394 190294 101450 190350
rect 101518 190294 101574 190350
rect 101642 190294 101698 190350
rect 101766 190294 101822 190350
rect 101394 190170 101450 190226
rect 101518 190170 101574 190226
rect 101642 190170 101698 190226
rect 101766 190170 101822 190226
rect 101394 190046 101450 190102
rect 101518 190046 101574 190102
rect 101642 190046 101698 190102
rect 101766 190046 101822 190102
rect 101394 189922 101450 189978
rect 101518 189922 101574 189978
rect 101642 189922 101698 189978
rect 101766 189922 101822 189978
rect 101394 172294 101450 172350
rect 101518 172294 101574 172350
rect 101642 172294 101698 172350
rect 101766 172294 101822 172350
rect 101394 172170 101450 172226
rect 101518 172170 101574 172226
rect 101642 172170 101698 172226
rect 101766 172170 101822 172226
rect 101394 172046 101450 172102
rect 101518 172046 101574 172102
rect 101642 172046 101698 172102
rect 101766 172046 101822 172102
rect 101394 171922 101450 171978
rect 101518 171922 101574 171978
rect 101642 171922 101698 171978
rect 101766 171922 101822 171978
rect 101394 154294 101450 154350
rect 101518 154294 101574 154350
rect 101642 154294 101698 154350
rect 101766 154294 101822 154350
rect 101394 154170 101450 154226
rect 101518 154170 101574 154226
rect 101642 154170 101698 154226
rect 101766 154170 101822 154226
rect 101394 154046 101450 154102
rect 101518 154046 101574 154102
rect 101642 154046 101698 154102
rect 101766 154046 101822 154102
rect 101394 153922 101450 153978
rect 101518 153922 101574 153978
rect 101642 153922 101698 153978
rect 101766 153922 101822 153978
rect 101394 136294 101450 136350
rect 101518 136294 101574 136350
rect 101642 136294 101698 136350
rect 101766 136294 101822 136350
rect 101394 136170 101450 136226
rect 101518 136170 101574 136226
rect 101642 136170 101698 136226
rect 101766 136170 101822 136226
rect 101394 136046 101450 136102
rect 101518 136046 101574 136102
rect 101642 136046 101698 136102
rect 101766 136046 101822 136102
rect 101394 135922 101450 135978
rect 101518 135922 101574 135978
rect 101642 135922 101698 135978
rect 101766 135922 101822 135978
rect 101394 118294 101450 118350
rect 101518 118294 101574 118350
rect 101642 118294 101698 118350
rect 101766 118294 101822 118350
rect 101394 118170 101450 118226
rect 101518 118170 101574 118226
rect 101642 118170 101698 118226
rect 101766 118170 101822 118226
rect 101394 118046 101450 118102
rect 101518 118046 101574 118102
rect 101642 118046 101698 118102
rect 101766 118046 101822 118102
rect 101394 117922 101450 117978
rect 101518 117922 101574 117978
rect 101642 117922 101698 117978
rect 101766 117922 101822 117978
rect 101394 100294 101450 100350
rect 101518 100294 101574 100350
rect 101642 100294 101698 100350
rect 101766 100294 101822 100350
rect 101394 100170 101450 100226
rect 101518 100170 101574 100226
rect 101642 100170 101698 100226
rect 101766 100170 101822 100226
rect 101394 100046 101450 100102
rect 101518 100046 101574 100102
rect 101642 100046 101698 100102
rect 101766 100046 101822 100102
rect 101394 99922 101450 99978
rect 101518 99922 101574 99978
rect 101642 99922 101698 99978
rect 101766 99922 101822 99978
rect 101394 82294 101450 82350
rect 101518 82294 101574 82350
rect 101642 82294 101698 82350
rect 101766 82294 101822 82350
rect 101394 82170 101450 82226
rect 101518 82170 101574 82226
rect 101642 82170 101698 82226
rect 101766 82170 101822 82226
rect 101394 82046 101450 82102
rect 101518 82046 101574 82102
rect 101642 82046 101698 82102
rect 101766 82046 101822 82102
rect 101394 81922 101450 81978
rect 101518 81922 101574 81978
rect 101642 81922 101698 81978
rect 101766 81922 101822 81978
rect 101394 64294 101450 64350
rect 101518 64294 101574 64350
rect 101642 64294 101698 64350
rect 101766 64294 101822 64350
rect 101394 64170 101450 64226
rect 101518 64170 101574 64226
rect 101642 64170 101698 64226
rect 101766 64170 101822 64226
rect 101394 64046 101450 64102
rect 101518 64046 101574 64102
rect 101642 64046 101698 64102
rect 101766 64046 101822 64102
rect 101394 63922 101450 63978
rect 101518 63922 101574 63978
rect 101642 63922 101698 63978
rect 101766 63922 101822 63978
rect 101394 46294 101450 46350
rect 101518 46294 101574 46350
rect 101642 46294 101698 46350
rect 101766 46294 101822 46350
rect 101394 46170 101450 46226
rect 101518 46170 101574 46226
rect 101642 46170 101698 46226
rect 101766 46170 101822 46226
rect 101394 46046 101450 46102
rect 101518 46046 101574 46102
rect 101642 46046 101698 46102
rect 101766 46046 101822 46102
rect 101394 45922 101450 45978
rect 101518 45922 101574 45978
rect 101642 45922 101698 45978
rect 101766 45922 101822 45978
rect 101394 28294 101450 28350
rect 101518 28294 101574 28350
rect 101642 28294 101698 28350
rect 101766 28294 101822 28350
rect 101394 28170 101450 28226
rect 101518 28170 101574 28226
rect 101642 28170 101698 28226
rect 101766 28170 101822 28226
rect 101394 28046 101450 28102
rect 101518 28046 101574 28102
rect 101642 28046 101698 28102
rect 101766 28046 101822 28102
rect 101394 27922 101450 27978
rect 101518 27922 101574 27978
rect 101642 27922 101698 27978
rect 101766 27922 101822 27978
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 110598 190294 110654 190350
rect 110722 190294 110778 190350
rect 110598 190170 110654 190226
rect 110722 190170 110778 190226
rect 110598 190046 110654 190102
rect 110722 190046 110778 190102
rect 110598 189922 110654 189978
rect 110722 189922 110778 189978
rect 110598 172294 110654 172350
rect 110722 172294 110778 172350
rect 110598 172170 110654 172226
rect 110722 172170 110778 172226
rect 110598 172046 110654 172102
rect 110722 172046 110778 172102
rect 110598 171922 110654 171978
rect 110722 171922 110778 171978
rect 114716 141002 114772 141058
rect 119308 142622 119364 142678
rect 119308 141902 119364 141958
rect 128394 274294 128450 274350
rect 128518 274294 128574 274350
rect 128642 274294 128698 274350
rect 128766 274294 128822 274350
rect 128394 274170 128450 274226
rect 128518 274170 128574 274226
rect 128642 274170 128698 274226
rect 128766 274170 128822 274226
rect 128394 274046 128450 274102
rect 128518 274046 128574 274102
rect 128642 274046 128698 274102
rect 128766 274046 128822 274102
rect 128394 273922 128450 273978
rect 128518 273922 128574 273978
rect 128642 273922 128698 273978
rect 128766 273922 128822 273978
rect 128394 256294 128450 256350
rect 128518 256294 128574 256350
rect 128642 256294 128698 256350
rect 128766 256294 128822 256350
rect 128394 256170 128450 256226
rect 128518 256170 128574 256226
rect 128642 256170 128698 256226
rect 128766 256170 128822 256226
rect 128394 256046 128450 256102
rect 128518 256046 128574 256102
rect 128642 256046 128698 256102
rect 128766 256046 128822 256102
rect 128394 255922 128450 255978
rect 128518 255922 128574 255978
rect 128642 255922 128698 255978
rect 128766 255922 128822 255978
rect 128394 238294 128450 238350
rect 128518 238294 128574 238350
rect 128642 238294 128698 238350
rect 128766 238294 128822 238350
rect 128394 238170 128450 238226
rect 128518 238170 128574 238226
rect 128642 238170 128698 238226
rect 128766 238170 128822 238226
rect 128394 238046 128450 238102
rect 128518 238046 128574 238102
rect 128642 238046 128698 238102
rect 128766 238046 128822 238102
rect 128394 237922 128450 237978
rect 128518 237922 128574 237978
rect 128642 237922 128698 237978
rect 128766 237922 128822 237978
rect 128394 220294 128450 220350
rect 128518 220294 128574 220350
rect 128642 220294 128698 220350
rect 128766 220294 128822 220350
rect 128394 220170 128450 220226
rect 128518 220170 128574 220226
rect 128642 220170 128698 220226
rect 128766 220170 128822 220226
rect 128394 220046 128450 220102
rect 128518 220046 128574 220102
rect 128642 220046 128698 220102
rect 128766 220046 128822 220102
rect 128394 219922 128450 219978
rect 128518 219922 128574 219978
rect 128642 219922 128698 219978
rect 128766 219922 128822 219978
rect 125958 202294 126014 202350
rect 126082 202294 126138 202350
rect 125958 202170 126014 202226
rect 126082 202170 126138 202226
rect 125958 202046 126014 202102
rect 126082 202046 126138 202102
rect 125958 201922 126014 201978
rect 126082 201922 126138 201978
rect 132114 298294 132170 298350
rect 132238 298294 132294 298350
rect 132362 298294 132418 298350
rect 132486 298294 132542 298350
rect 132114 298170 132170 298226
rect 132238 298170 132294 298226
rect 132362 298170 132418 298226
rect 132486 298170 132542 298226
rect 132114 298046 132170 298102
rect 132238 298046 132294 298102
rect 132362 298046 132418 298102
rect 132486 298046 132542 298102
rect 132114 297922 132170 297978
rect 132238 297922 132294 297978
rect 132362 297922 132418 297978
rect 132486 297922 132542 297978
rect 141318 298294 141374 298350
rect 141442 298294 141498 298350
rect 141318 298170 141374 298226
rect 141442 298170 141498 298226
rect 141318 298046 141374 298102
rect 141442 298046 141498 298102
rect 141318 297922 141374 297978
rect 141442 297922 141498 297978
rect 159114 292294 159170 292350
rect 159238 292294 159294 292350
rect 159362 292294 159418 292350
rect 159486 292294 159542 292350
rect 159114 292170 159170 292226
rect 159238 292170 159294 292226
rect 159362 292170 159418 292226
rect 159486 292170 159542 292226
rect 159114 292046 159170 292102
rect 159238 292046 159294 292102
rect 159362 292046 159418 292102
rect 159486 292046 159542 292102
rect 159114 291922 159170 291978
rect 159238 291922 159294 291978
rect 159362 291922 159418 291978
rect 159486 291922 159542 291978
rect 132114 280294 132170 280350
rect 132238 280294 132294 280350
rect 132362 280294 132418 280350
rect 132486 280294 132542 280350
rect 132114 280170 132170 280226
rect 132238 280170 132294 280226
rect 132362 280170 132418 280226
rect 132486 280170 132542 280226
rect 132114 280046 132170 280102
rect 132238 280046 132294 280102
rect 132362 280046 132418 280102
rect 132486 280046 132542 280102
rect 132114 279922 132170 279978
rect 132238 279922 132294 279978
rect 132362 279922 132418 279978
rect 132486 279922 132542 279978
rect 132114 262294 132170 262350
rect 132238 262294 132294 262350
rect 132362 262294 132418 262350
rect 132486 262294 132542 262350
rect 132114 262170 132170 262226
rect 132238 262170 132294 262226
rect 132362 262170 132418 262226
rect 132486 262170 132542 262226
rect 132114 262046 132170 262102
rect 132238 262046 132294 262102
rect 132362 262046 132418 262102
rect 132486 262046 132542 262102
rect 132114 261922 132170 261978
rect 132238 261922 132294 261978
rect 132362 261922 132418 261978
rect 132486 261922 132542 261978
rect 132114 244294 132170 244350
rect 132238 244294 132294 244350
rect 132362 244294 132418 244350
rect 132486 244294 132542 244350
rect 132114 244170 132170 244226
rect 132238 244170 132294 244226
rect 132362 244170 132418 244226
rect 132486 244170 132542 244226
rect 132114 244046 132170 244102
rect 132238 244046 132294 244102
rect 132362 244046 132418 244102
rect 132486 244046 132542 244102
rect 132114 243922 132170 243978
rect 132238 243922 132294 243978
rect 132362 243922 132418 243978
rect 132486 243922 132542 243978
rect 132114 226294 132170 226350
rect 132238 226294 132294 226350
rect 132362 226294 132418 226350
rect 132486 226294 132542 226350
rect 132114 226170 132170 226226
rect 132238 226170 132294 226226
rect 132362 226170 132418 226226
rect 132486 226170 132542 226226
rect 132114 226046 132170 226102
rect 132238 226046 132294 226102
rect 132362 226046 132418 226102
rect 132486 226046 132542 226102
rect 132114 225922 132170 225978
rect 132238 225922 132294 225978
rect 132362 225922 132418 225978
rect 132486 225922 132542 225978
rect 128394 202294 128450 202350
rect 128518 202294 128574 202350
rect 128642 202294 128698 202350
rect 128766 202294 128822 202350
rect 128394 202170 128450 202226
rect 128518 202170 128574 202226
rect 128642 202170 128698 202226
rect 128766 202170 128822 202226
rect 128394 202046 128450 202102
rect 128518 202046 128574 202102
rect 128642 202046 128698 202102
rect 128766 202046 128822 202102
rect 128394 201922 128450 201978
rect 128518 201922 128574 201978
rect 128642 201922 128698 201978
rect 128766 201922 128822 201978
rect 125958 184294 126014 184350
rect 126082 184294 126138 184350
rect 125958 184170 126014 184226
rect 126082 184170 126138 184226
rect 125958 184046 126014 184102
rect 126082 184046 126138 184102
rect 125958 183922 126014 183978
rect 126082 183922 126138 183978
rect 128394 184294 128450 184350
rect 128518 184294 128574 184350
rect 128642 184294 128698 184350
rect 128766 184294 128822 184350
rect 128394 184170 128450 184226
rect 128518 184170 128574 184226
rect 128642 184170 128698 184226
rect 128766 184170 128822 184226
rect 128394 184046 128450 184102
rect 128518 184046 128574 184102
rect 128642 184046 128698 184102
rect 128766 184046 128822 184102
rect 128394 183922 128450 183978
rect 128518 183922 128574 183978
rect 128642 183922 128698 183978
rect 128766 183922 128822 183978
rect 125958 166294 126014 166350
rect 126082 166294 126138 166350
rect 125958 166170 126014 166226
rect 126082 166170 126138 166226
rect 125958 166046 126014 166102
rect 126082 166046 126138 166102
rect 125958 165922 126014 165978
rect 126082 165922 126138 165978
rect 128394 166294 128450 166350
rect 128518 166294 128574 166350
rect 128642 166294 128698 166350
rect 128766 166294 128822 166350
rect 128394 166170 128450 166226
rect 128518 166170 128574 166226
rect 128642 166170 128698 166226
rect 128766 166170 128822 166226
rect 128394 166046 128450 166102
rect 128518 166046 128574 166102
rect 128642 166046 128698 166102
rect 128766 166046 128822 166102
rect 128394 165922 128450 165978
rect 128518 165922 128574 165978
rect 128642 165922 128698 165978
rect 128766 165922 128822 165978
rect 128394 148294 128450 148350
rect 128518 148294 128574 148350
rect 128642 148294 128698 148350
rect 128766 148294 128822 148350
rect 128394 148170 128450 148226
rect 128518 148170 128574 148226
rect 128642 148170 128698 148226
rect 128766 148170 128822 148226
rect 128394 148046 128450 148102
rect 128518 148046 128574 148102
rect 128642 148046 128698 148102
rect 128766 148046 128822 148102
rect 128394 147922 128450 147978
rect 128518 147922 128574 147978
rect 128642 147922 128698 147978
rect 128766 147922 128822 147978
rect 128394 130294 128450 130350
rect 128518 130294 128574 130350
rect 128642 130294 128698 130350
rect 128766 130294 128822 130350
rect 128394 130170 128450 130226
rect 128518 130170 128574 130226
rect 128642 130170 128698 130226
rect 128766 130170 128822 130226
rect 128394 130046 128450 130102
rect 128518 130046 128574 130102
rect 128642 130046 128698 130102
rect 128766 130046 128822 130102
rect 128394 129922 128450 129978
rect 128518 129922 128574 129978
rect 128642 129922 128698 129978
rect 128766 129922 128822 129978
rect 128394 112294 128450 112350
rect 128518 112294 128574 112350
rect 128642 112294 128698 112350
rect 128766 112294 128822 112350
rect 128394 112170 128450 112226
rect 128518 112170 128574 112226
rect 128642 112170 128698 112226
rect 128766 112170 128822 112226
rect 128394 112046 128450 112102
rect 128518 112046 128574 112102
rect 128642 112046 128698 112102
rect 128766 112046 128822 112102
rect 128394 111922 128450 111978
rect 128518 111922 128574 111978
rect 128642 111922 128698 111978
rect 128766 111922 128822 111978
rect 128394 94294 128450 94350
rect 128518 94294 128574 94350
rect 128642 94294 128698 94350
rect 128766 94294 128822 94350
rect 128394 94170 128450 94226
rect 128518 94170 128574 94226
rect 128642 94170 128698 94226
rect 128766 94170 128822 94226
rect 128394 94046 128450 94102
rect 128518 94046 128574 94102
rect 128642 94046 128698 94102
rect 128766 94046 128822 94102
rect 128394 93922 128450 93978
rect 128518 93922 128574 93978
rect 128642 93922 128698 93978
rect 128766 93922 128822 93978
rect 128394 76294 128450 76350
rect 128518 76294 128574 76350
rect 128642 76294 128698 76350
rect 128766 76294 128822 76350
rect 128394 76170 128450 76226
rect 128518 76170 128574 76226
rect 128642 76170 128698 76226
rect 128766 76170 128822 76226
rect 128394 76046 128450 76102
rect 128518 76046 128574 76102
rect 128642 76046 128698 76102
rect 128766 76046 128822 76102
rect 128394 75922 128450 75978
rect 128518 75922 128574 75978
rect 128642 75922 128698 75978
rect 128766 75922 128822 75978
rect 128394 58294 128450 58350
rect 128518 58294 128574 58350
rect 128642 58294 128698 58350
rect 128766 58294 128822 58350
rect 128394 58170 128450 58226
rect 128518 58170 128574 58226
rect 128642 58170 128698 58226
rect 128766 58170 128822 58226
rect 128394 58046 128450 58102
rect 128518 58046 128574 58102
rect 128642 58046 128698 58102
rect 128766 58046 128822 58102
rect 128394 57922 128450 57978
rect 128518 57922 128574 57978
rect 128642 57922 128698 57978
rect 128766 57922 128822 57978
rect 128394 40294 128450 40350
rect 128518 40294 128574 40350
rect 128642 40294 128698 40350
rect 128766 40294 128822 40350
rect 128394 40170 128450 40226
rect 128518 40170 128574 40226
rect 128642 40170 128698 40226
rect 128766 40170 128822 40226
rect 128394 40046 128450 40102
rect 128518 40046 128574 40102
rect 128642 40046 128698 40102
rect 128766 40046 128822 40102
rect 128394 39922 128450 39978
rect 128518 39922 128574 39978
rect 128642 39922 128698 39978
rect 128766 39922 128822 39978
rect 128394 22294 128450 22350
rect 128518 22294 128574 22350
rect 128642 22294 128698 22350
rect 128766 22294 128822 22350
rect 128394 22170 128450 22226
rect 128518 22170 128574 22226
rect 128642 22170 128698 22226
rect 128766 22170 128822 22226
rect 128394 22046 128450 22102
rect 128518 22046 128574 22102
rect 128642 22046 128698 22102
rect 128766 22046 128822 22102
rect 128394 21922 128450 21978
rect 128518 21922 128574 21978
rect 128642 21922 128698 21978
rect 128766 21922 128822 21978
rect 132114 208294 132170 208350
rect 132238 208294 132294 208350
rect 132362 208294 132418 208350
rect 132486 208294 132542 208350
rect 132114 208170 132170 208226
rect 132238 208170 132294 208226
rect 132362 208170 132418 208226
rect 132486 208170 132542 208226
rect 132114 208046 132170 208102
rect 132238 208046 132294 208102
rect 132362 208046 132418 208102
rect 132486 208046 132542 208102
rect 132114 207922 132170 207978
rect 132238 207922 132294 207978
rect 132362 207922 132418 207978
rect 132486 207922 132542 207978
rect 132114 190294 132170 190350
rect 132238 190294 132294 190350
rect 132362 190294 132418 190350
rect 132486 190294 132542 190350
rect 132114 190170 132170 190226
rect 132238 190170 132294 190226
rect 132362 190170 132418 190226
rect 132486 190170 132542 190226
rect 132114 190046 132170 190102
rect 132238 190046 132294 190102
rect 132362 190046 132418 190102
rect 132486 190046 132542 190102
rect 132114 189922 132170 189978
rect 132238 189922 132294 189978
rect 132362 189922 132418 189978
rect 132486 189922 132542 189978
rect 132114 172294 132170 172350
rect 132238 172294 132294 172350
rect 132362 172294 132418 172350
rect 132486 172294 132542 172350
rect 132114 172170 132170 172226
rect 132238 172170 132294 172226
rect 132362 172170 132418 172226
rect 132486 172170 132542 172226
rect 132114 172046 132170 172102
rect 132238 172046 132294 172102
rect 132362 172046 132418 172102
rect 132486 172046 132542 172102
rect 132114 171922 132170 171978
rect 132238 171922 132294 171978
rect 132362 171922 132418 171978
rect 132486 171922 132542 171978
rect 132114 154294 132170 154350
rect 132238 154294 132294 154350
rect 132362 154294 132418 154350
rect 132486 154294 132542 154350
rect 132114 154170 132170 154226
rect 132238 154170 132294 154226
rect 132362 154170 132418 154226
rect 132486 154170 132542 154226
rect 132114 154046 132170 154102
rect 132238 154046 132294 154102
rect 132362 154046 132418 154102
rect 132486 154046 132542 154102
rect 132114 153922 132170 153978
rect 132238 153922 132294 153978
rect 132362 153922 132418 153978
rect 132486 153922 132542 153978
rect 130956 142268 131012 142318
rect 130956 142262 131012 142268
rect 132114 136294 132170 136350
rect 132238 136294 132294 136350
rect 132362 136294 132418 136350
rect 132486 136294 132542 136350
rect 132114 136170 132170 136226
rect 132238 136170 132294 136226
rect 132362 136170 132418 136226
rect 132486 136170 132542 136226
rect 132114 136046 132170 136102
rect 132238 136046 132294 136102
rect 132362 136046 132418 136102
rect 132486 136046 132542 136102
rect 132114 135922 132170 135978
rect 132238 135922 132294 135978
rect 132362 135922 132418 135978
rect 132486 135922 132542 135978
rect 132114 118294 132170 118350
rect 132238 118294 132294 118350
rect 132362 118294 132418 118350
rect 132486 118294 132542 118350
rect 132114 118170 132170 118226
rect 132238 118170 132294 118226
rect 132362 118170 132418 118226
rect 132486 118170 132542 118226
rect 132114 118046 132170 118102
rect 132238 118046 132294 118102
rect 132362 118046 132418 118102
rect 132486 118046 132542 118102
rect 132114 117922 132170 117978
rect 132238 117922 132294 117978
rect 132362 117922 132418 117978
rect 132486 117922 132542 117978
rect 132114 100294 132170 100350
rect 132238 100294 132294 100350
rect 132362 100294 132418 100350
rect 132486 100294 132542 100350
rect 132114 100170 132170 100226
rect 132238 100170 132294 100226
rect 132362 100170 132418 100226
rect 132486 100170 132542 100226
rect 132114 100046 132170 100102
rect 132238 100046 132294 100102
rect 132362 100046 132418 100102
rect 132486 100046 132542 100102
rect 132114 99922 132170 99978
rect 132238 99922 132294 99978
rect 132362 99922 132418 99978
rect 132486 99922 132542 99978
rect 132114 82294 132170 82350
rect 132238 82294 132294 82350
rect 132362 82294 132418 82350
rect 132486 82294 132542 82350
rect 132114 82170 132170 82226
rect 132238 82170 132294 82226
rect 132362 82170 132418 82226
rect 132486 82170 132542 82226
rect 132114 82046 132170 82102
rect 132238 82046 132294 82102
rect 132362 82046 132418 82102
rect 132486 82046 132542 82102
rect 132114 81922 132170 81978
rect 132238 81922 132294 81978
rect 132362 81922 132418 81978
rect 132486 81922 132542 81978
rect 132114 64294 132170 64350
rect 132238 64294 132294 64350
rect 132362 64294 132418 64350
rect 132486 64294 132542 64350
rect 132114 64170 132170 64226
rect 132238 64170 132294 64226
rect 132362 64170 132418 64226
rect 132486 64170 132542 64226
rect 132114 64046 132170 64102
rect 132238 64046 132294 64102
rect 132362 64046 132418 64102
rect 132486 64046 132542 64102
rect 132114 63922 132170 63978
rect 132238 63922 132294 63978
rect 132362 63922 132418 63978
rect 132486 63922 132542 63978
rect 132114 46294 132170 46350
rect 132238 46294 132294 46350
rect 132362 46294 132418 46350
rect 132486 46294 132542 46350
rect 132114 46170 132170 46226
rect 132238 46170 132294 46226
rect 132362 46170 132418 46226
rect 132486 46170 132542 46226
rect 132114 46046 132170 46102
rect 132238 46046 132294 46102
rect 132362 46046 132418 46102
rect 132486 46046 132542 46102
rect 132114 45922 132170 45978
rect 132238 45922 132294 45978
rect 132362 45922 132418 45978
rect 132486 45922 132542 45978
rect 132114 28294 132170 28350
rect 132238 28294 132294 28350
rect 132362 28294 132418 28350
rect 132486 28294 132542 28350
rect 132114 28170 132170 28226
rect 132238 28170 132294 28226
rect 132362 28170 132418 28226
rect 132486 28170 132542 28226
rect 132114 28046 132170 28102
rect 132238 28046 132294 28102
rect 132362 28046 132418 28102
rect 132486 28046 132542 28102
rect 132114 27922 132170 27978
rect 132238 27922 132294 27978
rect 132362 27922 132418 27978
rect 132486 27922 132542 27978
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 141318 190294 141374 190350
rect 141442 190294 141498 190350
rect 141318 190170 141374 190226
rect 141442 190170 141498 190226
rect 141318 190046 141374 190102
rect 141442 190046 141498 190102
rect 141318 189922 141374 189978
rect 141442 189922 141498 189978
rect 141318 172294 141374 172350
rect 141442 172294 141498 172350
rect 141318 172170 141374 172226
rect 141442 172170 141498 172226
rect 141318 172046 141374 172102
rect 141442 172046 141498 172102
rect 141318 171922 141374 171978
rect 141442 171922 141498 171978
rect 144732 142622 144788 142678
rect 145404 140822 145460 140878
rect 145812 130294 145868 130350
rect 145936 130294 145992 130350
rect 146060 130294 146116 130350
rect 146184 130294 146240 130350
rect 145812 130170 145868 130226
rect 145936 130170 145992 130226
rect 146060 130170 146116 130226
rect 146184 130170 146240 130226
rect 145812 130046 145868 130102
rect 145936 130046 145992 130102
rect 146060 130046 146116 130102
rect 146184 130046 146240 130102
rect 145812 129922 145868 129978
rect 145936 129922 145992 129978
rect 146060 129922 146116 129978
rect 146184 129922 146240 129978
rect 146612 118294 146668 118350
rect 146736 118294 146792 118350
rect 146860 118294 146916 118350
rect 146984 118294 147040 118350
rect 146612 118170 146668 118226
rect 146736 118170 146792 118226
rect 146860 118170 146916 118226
rect 146984 118170 147040 118226
rect 146612 118046 146668 118102
rect 146736 118046 146792 118102
rect 146860 118046 146916 118102
rect 146984 118046 147040 118102
rect 146612 117922 146668 117978
rect 146736 117922 146792 117978
rect 146860 117922 146916 117978
rect 146984 117922 147040 117978
rect 145812 112294 145868 112350
rect 145936 112294 145992 112350
rect 146060 112294 146116 112350
rect 146184 112294 146240 112350
rect 145812 112170 145868 112226
rect 145936 112170 145992 112226
rect 146060 112170 146116 112226
rect 146184 112170 146240 112226
rect 145812 112046 145868 112102
rect 145936 112046 145992 112102
rect 146060 112046 146116 112102
rect 146184 112046 146240 112102
rect 145812 111922 145868 111978
rect 145936 111922 145992 111978
rect 146060 111922 146116 111978
rect 146184 111922 146240 111978
rect 146612 100294 146668 100350
rect 146736 100294 146792 100350
rect 146860 100294 146916 100350
rect 146984 100294 147040 100350
rect 146612 100170 146668 100226
rect 146736 100170 146792 100226
rect 146860 100170 146916 100226
rect 146984 100170 147040 100226
rect 146612 100046 146668 100102
rect 146736 100046 146792 100102
rect 146860 100046 146916 100102
rect 146984 100046 147040 100102
rect 146612 99922 146668 99978
rect 146736 99922 146792 99978
rect 146860 99922 146916 99978
rect 146984 99922 147040 99978
rect 145812 94294 145868 94350
rect 145936 94294 145992 94350
rect 146060 94294 146116 94350
rect 146184 94294 146240 94350
rect 145812 94170 145868 94226
rect 145936 94170 145992 94226
rect 146060 94170 146116 94226
rect 146184 94170 146240 94226
rect 145812 94046 145868 94102
rect 145936 94046 145992 94102
rect 146060 94046 146116 94102
rect 146184 94046 146240 94102
rect 145812 93922 145868 93978
rect 145936 93922 145992 93978
rect 146060 93922 146116 93978
rect 146184 93922 146240 93978
rect 146612 82294 146668 82350
rect 146736 82294 146792 82350
rect 146860 82294 146916 82350
rect 146984 82294 147040 82350
rect 146612 82170 146668 82226
rect 146736 82170 146792 82226
rect 146860 82170 146916 82226
rect 146984 82170 147040 82226
rect 146612 82046 146668 82102
rect 146736 82046 146792 82102
rect 146860 82046 146916 82102
rect 146984 82046 147040 82102
rect 146612 81922 146668 81978
rect 146736 81922 146792 81978
rect 146860 81922 146916 81978
rect 146984 81922 147040 81978
rect 145812 76294 145868 76350
rect 145936 76294 145992 76350
rect 146060 76294 146116 76350
rect 146184 76294 146240 76350
rect 145812 76170 145868 76226
rect 145936 76170 145992 76226
rect 146060 76170 146116 76226
rect 146184 76170 146240 76226
rect 145812 76046 145868 76102
rect 145936 76046 145992 76102
rect 146060 76046 146116 76102
rect 146184 76046 146240 76102
rect 145812 75922 145868 75978
rect 145936 75922 145992 75978
rect 146060 75922 146116 75978
rect 146184 75922 146240 75978
rect 146612 64294 146668 64350
rect 146736 64294 146792 64350
rect 146860 64294 146916 64350
rect 146984 64294 147040 64350
rect 146612 64170 146668 64226
rect 146736 64170 146792 64226
rect 146860 64170 146916 64226
rect 146984 64170 147040 64226
rect 146612 64046 146668 64102
rect 146736 64046 146792 64102
rect 146860 64046 146916 64102
rect 146984 64046 147040 64102
rect 146612 63922 146668 63978
rect 146736 63922 146792 63978
rect 146860 63922 146916 63978
rect 146984 63922 147040 63978
rect 145812 58294 145868 58350
rect 145936 58294 145992 58350
rect 146060 58294 146116 58350
rect 146184 58294 146240 58350
rect 145812 58170 145868 58226
rect 145936 58170 145992 58226
rect 146060 58170 146116 58226
rect 146184 58170 146240 58226
rect 145812 58046 145868 58102
rect 145936 58046 145992 58102
rect 146060 58046 146116 58102
rect 146184 58046 146240 58102
rect 145812 57922 145868 57978
rect 145936 57922 145992 57978
rect 146060 57922 146116 57978
rect 146184 57922 146240 57978
rect 146612 46294 146668 46350
rect 146736 46294 146792 46350
rect 146860 46294 146916 46350
rect 146984 46294 147040 46350
rect 146612 46170 146668 46226
rect 146736 46170 146792 46226
rect 146860 46170 146916 46226
rect 146984 46170 147040 46226
rect 146612 46046 146668 46102
rect 146736 46046 146792 46102
rect 146860 46046 146916 46102
rect 146984 46046 147040 46102
rect 146612 45922 146668 45978
rect 146736 45922 146792 45978
rect 146860 45922 146916 45978
rect 146984 45922 147040 45978
rect 152124 167282 152180 167338
rect 162834 298294 162890 298350
rect 162958 298294 163014 298350
rect 163082 298294 163138 298350
rect 163206 298294 163262 298350
rect 162834 298170 162890 298226
rect 162958 298170 163014 298226
rect 163082 298170 163138 298226
rect 163206 298170 163262 298226
rect 162834 298046 162890 298102
rect 162958 298046 163014 298102
rect 163082 298046 163138 298102
rect 163206 298046 163262 298102
rect 162834 297922 162890 297978
rect 162958 297922 163014 297978
rect 163082 297922 163138 297978
rect 163206 297922 163262 297978
rect 159114 274294 159170 274350
rect 159238 274294 159294 274350
rect 159362 274294 159418 274350
rect 159486 274294 159542 274350
rect 159114 274170 159170 274226
rect 159238 274170 159294 274226
rect 159362 274170 159418 274226
rect 159486 274170 159542 274226
rect 159114 274046 159170 274102
rect 159238 274046 159294 274102
rect 159362 274046 159418 274102
rect 159486 274046 159542 274102
rect 159114 273922 159170 273978
rect 159238 273922 159294 273978
rect 159362 273922 159418 273978
rect 159486 273922 159542 273978
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 156678 202294 156734 202350
rect 156802 202294 156858 202350
rect 156678 202170 156734 202226
rect 156802 202170 156858 202226
rect 156678 202046 156734 202102
rect 156802 202046 156858 202102
rect 156678 201922 156734 201978
rect 156802 201922 156858 201978
rect 159114 202294 159170 202350
rect 159238 202294 159294 202350
rect 159362 202294 159418 202350
rect 159486 202294 159542 202350
rect 159114 202170 159170 202226
rect 159238 202170 159294 202226
rect 159362 202170 159418 202226
rect 159486 202170 159542 202226
rect 159114 202046 159170 202102
rect 159238 202046 159294 202102
rect 159362 202046 159418 202102
rect 159486 202046 159542 202102
rect 159114 201922 159170 201978
rect 159238 201922 159294 201978
rect 159362 201922 159418 201978
rect 159486 201922 159542 201978
rect 156678 184294 156734 184350
rect 156802 184294 156858 184350
rect 156678 184170 156734 184226
rect 156802 184170 156858 184226
rect 156678 184046 156734 184102
rect 156802 184046 156858 184102
rect 156678 183922 156734 183978
rect 156802 183922 156858 183978
rect 159114 184294 159170 184350
rect 159238 184294 159294 184350
rect 159362 184294 159418 184350
rect 159486 184294 159542 184350
rect 159114 184170 159170 184226
rect 159238 184170 159294 184226
rect 159362 184170 159418 184226
rect 159486 184170 159542 184226
rect 159114 184046 159170 184102
rect 159238 184046 159294 184102
rect 159362 184046 159418 184102
rect 159486 184046 159542 184102
rect 159114 183922 159170 183978
rect 159238 183922 159294 183978
rect 159362 183922 159418 183978
rect 159486 183922 159542 183978
rect 157052 168722 157108 168778
rect 156678 166294 156734 166350
rect 156802 166294 156858 166350
rect 156678 166170 156734 166226
rect 156802 166170 156858 166226
rect 156678 166046 156734 166102
rect 156802 166046 156858 166102
rect 156678 165922 156734 165978
rect 156802 165922 156858 165978
rect 137228 4922 137284 4978
rect 155484 4922 155540 4978
rect 159114 166294 159170 166350
rect 159238 166294 159294 166350
rect 159362 166294 159418 166350
rect 159486 166294 159542 166350
rect 159114 166170 159170 166226
rect 159238 166170 159294 166226
rect 159362 166170 159418 166226
rect 159486 166170 159542 166226
rect 159114 166046 159170 166102
rect 159238 166046 159294 166102
rect 159362 166046 159418 166102
rect 159486 166046 159542 166102
rect 159114 165922 159170 165978
rect 159238 165922 159294 165978
rect 159362 165922 159418 165978
rect 159486 165922 159542 165978
rect 159114 148294 159170 148350
rect 159238 148294 159294 148350
rect 159362 148294 159418 148350
rect 159486 148294 159542 148350
rect 159114 148170 159170 148226
rect 159238 148170 159294 148226
rect 159362 148170 159418 148226
rect 159486 148170 159542 148226
rect 159114 148046 159170 148102
rect 159238 148046 159294 148102
rect 159362 148046 159418 148102
rect 159486 148046 159542 148102
rect 159114 147922 159170 147978
rect 159238 147922 159294 147978
rect 159362 147922 159418 147978
rect 159486 147922 159542 147978
rect 159114 130294 159170 130350
rect 159238 130294 159294 130350
rect 159362 130294 159418 130350
rect 159486 130294 159542 130350
rect 159114 130170 159170 130226
rect 159238 130170 159294 130226
rect 159362 130170 159418 130226
rect 159486 130170 159542 130226
rect 159114 130046 159170 130102
rect 159238 130046 159294 130102
rect 159362 130046 159418 130102
rect 159486 130046 159542 130102
rect 159114 129922 159170 129978
rect 159238 129922 159294 129978
rect 159362 129922 159418 129978
rect 159486 129922 159542 129978
rect 159114 112294 159170 112350
rect 159238 112294 159294 112350
rect 159362 112294 159418 112350
rect 159486 112294 159542 112350
rect 159114 112170 159170 112226
rect 159238 112170 159294 112226
rect 159362 112170 159418 112226
rect 159486 112170 159542 112226
rect 159114 112046 159170 112102
rect 159238 112046 159294 112102
rect 159362 112046 159418 112102
rect 159486 112046 159542 112102
rect 159114 111922 159170 111978
rect 159238 111922 159294 111978
rect 159362 111922 159418 111978
rect 159486 111922 159542 111978
rect 159114 94294 159170 94350
rect 159238 94294 159294 94350
rect 159362 94294 159418 94350
rect 159486 94294 159542 94350
rect 159114 94170 159170 94226
rect 159238 94170 159294 94226
rect 159362 94170 159418 94226
rect 159486 94170 159542 94226
rect 159114 94046 159170 94102
rect 159238 94046 159294 94102
rect 159362 94046 159418 94102
rect 159486 94046 159542 94102
rect 159114 93922 159170 93978
rect 159238 93922 159294 93978
rect 159362 93922 159418 93978
rect 159486 93922 159542 93978
rect 159114 76294 159170 76350
rect 159238 76294 159294 76350
rect 159362 76294 159418 76350
rect 159486 76294 159542 76350
rect 159114 76170 159170 76226
rect 159238 76170 159294 76226
rect 159362 76170 159418 76226
rect 159486 76170 159542 76226
rect 159114 76046 159170 76102
rect 159238 76046 159294 76102
rect 159362 76046 159418 76102
rect 159486 76046 159542 76102
rect 159114 75922 159170 75978
rect 159238 75922 159294 75978
rect 159362 75922 159418 75978
rect 159486 75922 159542 75978
rect 159114 58294 159170 58350
rect 159238 58294 159294 58350
rect 159362 58294 159418 58350
rect 159486 58294 159542 58350
rect 159114 58170 159170 58226
rect 159238 58170 159294 58226
rect 159362 58170 159418 58226
rect 159486 58170 159542 58226
rect 159114 58046 159170 58102
rect 159238 58046 159294 58102
rect 159362 58046 159418 58102
rect 159486 58046 159542 58102
rect 159114 57922 159170 57978
rect 159238 57922 159294 57978
rect 159362 57922 159418 57978
rect 159486 57922 159542 57978
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 172038 298294 172094 298350
rect 172162 298294 172218 298350
rect 172038 298170 172094 298226
rect 172162 298170 172218 298226
rect 172038 298046 172094 298102
rect 172162 298046 172218 298102
rect 172038 297922 172094 297978
rect 172162 297922 172218 297978
rect 189834 292294 189890 292350
rect 189958 292294 190014 292350
rect 190082 292294 190138 292350
rect 190206 292294 190262 292350
rect 189834 292170 189890 292226
rect 189958 292170 190014 292226
rect 190082 292170 190138 292226
rect 190206 292170 190262 292226
rect 189834 292046 189890 292102
rect 189958 292046 190014 292102
rect 190082 292046 190138 292102
rect 190206 292046 190262 292102
rect 189834 291922 189890 291978
rect 189958 291922 190014 291978
rect 190082 291922 190138 291978
rect 190206 291922 190262 291978
rect 162834 280294 162890 280350
rect 162958 280294 163014 280350
rect 163082 280294 163138 280350
rect 163206 280294 163262 280350
rect 162834 280170 162890 280226
rect 162958 280170 163014 280226
rect 163082 280170 163138 280226
rect 163206 280170 163262 280226
rect 162834 280046 162890 280102
rect 162958 280046 163014 280102
rect 163082 280046 163138 280102
rect 163206 280046 163262 280102
rect 162834 279922 162890 279978
rect 162958 279922 163014 279978
rect 163082 279922 163138 279978
rect 163206 279922 163262 279978
rect 162834 262294 162890 262350
rect 162958 262294 163014 262350
rect 163082 262294 163138 262350
rect 163206 262294 163262 262350
rect 162834 262170 162890 262226
rect 162958 262170 163014 262226
rect 163082 262170 163138 262226
rect 163206 262170 163262 262226
rect 162834 262046 162890 262102
rect 162958 262046 163014 262102
rect 163082 262046 163138 262102
rect 163206 262046 163262 262102
rect 162834 261922 162890 261978
rect 162958 261922 163014 261978
rect 163082 261922 163138 261978
rect 163206 261922 163262 261978
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 162834 208294 162890 208350
rect 162958 208294 163014 208350
rect 163082 208294 163138 208350
rect 163206 208294 163262 208350
rect 162834 208170 162890 208226
rect 162958 208170 163014 208226
rect 163082 208170 163138 208226
rect 163206 208170 163262 208226
rect 162834 208046 162890 208102
rect 162958 208046 163014 208102
rect 163082 208046 163138 208102
rect 163206 208046 163262 208102
rect 162834 207922 162890 207978
rect 162958 207922 163014 207978
rect 163082 207922 163138 207978
rect 163206 207922 163262 207978
rect 162834 190294 162890 190350
rect 162958 190294 163014 190350
rect 163082 190294 163138 190350
rect 163206 190294 163262 190350
rect 162834 190170 162890 190226
rect 162958 190170 163014 190226
rect 163082 190170 163138 190226
rect 163206 190170 163262 190226
rect 162834 190046 162890 190102
rect 162958 190046 163014 190102
rect 163082 190046 163138 190102
rect 163206 190046 163262 190102
rect 162834 189922 162890 189978
rect 162958 189922 163014 189978
rect 163082 189922 163138 189978
rect 163206 189922 163262 189978
rect 160412 173762 160468 173818
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 162834 172294 162890 172350
rect 162958 172294 163014 172350
rect 163082 172294 163138 172350
rect 163206 172294 163262 172350
rect 162834 172170 162890 172226
rect 162958 172170 163014 172226
rect 163082 172170 163138 172226
rect 163206 172170 163262 172226
rect 162834 172046 162890 172102
rect 162958 172046 163014 172102
rect 163082 172046 163138 172102
rect 163206 172046 163262 172102
rect 162834 171922 162890 171978
rect 162958 171922 163014 171978
rect 163082 171922 163138 171978
rect 163206 171922 163262 171978
rect 162834 154294 162890 154350
rect 162958 154294 163014 154350
rect 163082 154294 163138 154350
rect 163206 154294 163262 154350
rect 162834 154170 162890 154226
rect 162958 154170 163014 154226
rect 163082 154170 163138 154226
rect 163206 154170 163262 154226
rect 162834 154046 162890 154102
rect 162958 154046 163014 154102
rect 163082 154046 163138 154102
rect 163206 154046 163262 154102
rect 162834 153922 162890 153978
rect 162958 153922 163014 153978
rect 163082 153922 163138 153978
rect 163206 153922 163262 153978
rect 167916 170522 167972 170578
rect 164444 142082 164500 142138
rect 162834 136294 162890 136350
rect 162958 136294 163014 136350
rect 163082 136294 163138 136350
rect 163206 136294 163262 136350
rect 162834 136170 162890 136226
rect 162958 136170 163014 136226
rect 163082 136170 163138 136226
rect 163206 136170 163262 136226
rect 162834 136046 162890 136102
rect 162958 136046 163014 136102
rect 163082 136046 163138 136102
rect 163206 136046 163262 136102
rect 162834 135922 162890 135978
rect 162958 135922 163014 135978
rect 163082 135922 163138 135978
rect 163206 135922 163262 135978
rect 161130 130294 161186 130350
rect 161254 130294 161310 130350
rect 161378 130294 161434 130350
rect 161502 130294 161558 130350
rect 161130 130170 161186 130226
rect 161254 130170 161310 130226
rect 161378 130170 161434 130226
rect 161502 130170 161558 130226
rect 161130 130046 161186 130102
rect 161254 130046 161310 130102
rect 161378 130046 161434 130102
rect 161502 130046 161558 130102
rect 161130 129922 161186 129978
rect 161254 129922 161310 129978
rect 161378 129922 161434 129978
rect 161502 129922 161558 129978
rect 161930 118294 161986 118350
rect 162054 118294 162110 118350
rect 162178 118294 162234 118350
rect 162302 118294 162358 118350
rect 161930 118170 161986 118226
rect 162054 118170 162110 118226
rect 162178 118170 162234 118226
rect 162302 118170 162358 118226
rect 161930 118046 161986 118102
rect 162054 118046 162110 118102
rect 162178 118046 162234 118102
rect 162302 118046 162358 118102
rect 161930 117922 161986 117978
rect 162054 117922 162110 117978
rect 162178 117922 162234 117978
rect 162302 117922 162358 117978
rect 162834 118294 162890 118350
rect 162958 118294 163014 118350
rect 163082 118294 163138 118350
rect 163206 118294 163262 118350
rect 162834 118170 162890 118226
rect 162958 118170 163014 118226
rect 163082 118170 163138 118226
rect 163206 118170 163262 118226
rect 162834 118046 162890 118102
rect 162958 118046 163014 118102
rect 163082 118046 163138 118102
rect 163206 118046 163262 118102
rect 162834 117922 162890 117978
rect 162958 117922 163014 117978
rect 163082 117922 163138 117978
rect 163206 117922 163262 117978
rect 161130 112294 161186 112350
rect 161254 112294 161310 112350
rect 161378 112294 161434 112350
rect 161502 112294 161558 112350
rect 161130 112170 161186 112226
rect 161254 112170 161310 112226
rect 161378 112170 161434 112226
rect 161502 112170 161558 112226
rect 161130 112046 161186 112102
rect 161254 112046 161310 112102
rect 161378 112046 161434 112102
rect 161502 112046 161558 112102
rect 161130 111922 161186 111978
rect 161254 111922 161310 111978
rect 161378 111922 161434 111978
rect 161502 111922 161558 111978
rect 161930 100294 161986 100350
rect 162054 100294 162110 100350
rect 162178 100294 162234 100350
rect 162302 100294 162358 100350
rect 161930 100170 161986 100226
rect 162054 100170 162110 100226
rect 162178 100170 162234 100226
rect 162302 100170 162358 100226
rect 161930 100046 161986 100102
rect 162054 100046 162110 100102
rect 162178 100046 162234 100102
rect 162302 100046 162358 100102
rect 161930 99922 161986 99978
rect 162054 99922 162110 99978
rect 162178 99922 162234 99978
rect 162302 99922 162358 99978
rect 162834 100294 162890 100350
rect 162958 100294 163014 100350
rect 163082 100294 163138 100350
rect 163206 100294 163262 100350
rect 162834 100170 162890 100226
rect 162958 100170 163014 100226
rect 163082 100170 163138 100226
rect 163206 100170 163262 100226
rect 162834 100046 162890 100102
rect 162958 100046 163014 100102
rect 163082 100046 163138 100102
rect 163206 100046 163262 100102
rect 162834 99922 162890 99978
rect 162958 99922 163014 99978
rect 163082 99922 163138 99978
rect 163206 99922 163262 99978
rect 161130 94294 161186 94350
rect 161254 94294 161310 94350
rect 161378 94294 161434 94350
rect 161502 94294 161558 94350
rect 161130 94170 161186 94226
rect 161254 94170 161310 94226
rect 161378 94170 161434 94226
rect 161502 94170 161558 94226
rect 161130 94046 161186 94102
rect 161254 94046 161310 94102
rect 161378 94046 161434 94102
rect 161502 94046 161558 94102
rect 161130 93922 161186 93978
rect 161254 93922 161310 93978
rect 161378 93922 161434 93978
rect 161502 93922 161558 93978
rect 161930 82294 161986 82350
rect 162054 82294 162110 82350
rect 162178 82294 162234 82350
rect 162302 82294 162358 82350
rect 161930 82170 161986 82226
rect 162054 82170 162110 82226
rect 162178 82170 162234 82226
rect 162302 82170 162358 82226
rect 161930 82046 161986 82102
rect 162054 82046 162110 82102
rect 162178 82046 162234 82102
rect 162302 82046 162358 82102
rect 161930 81922 161986 81978
rect 162054 81922 162110 81978
rect 162178 81922 162234 81978
rect 162302 81922 162358 81978
rect 162834 82294 162890 82350
rect 162958 82294 163014 82350
rect 163082 82294 163138 82350
rect 163206 82294 163262 82350
rect 162834 82170 162890 82226
rect 162958 82170 163014 82226
rect 163082 82170 163138 82226
rect 163206 82170 163262 82226
rect 162834 82046 162890 82102
rect 162958 82046 163014 82102
rect 163082 82046 163138 82102
rect 163206 82046 163262 82102
rect 162834 81922 162890 81978
rect 162958 81922 163014 81978
rect 163082 81922 163138 81978
rect 163206 81922 163262 81978
rect 161130 76294 161186 76350
rect 161254 76294 161310 76350
rect 161378 76294 161434 76350
rect 161502 76294 161558 76350
rect 161130 76170 161186 76226
rect 161254 76170 161310 76226
rect 161378 76170 161434 76226
rect 161502 76170 161558 76226
rect 161130 76046 161186 76102
rect 161254 76046 161310 76102
rect 161378 76046 161434 76102
rect 161502 76046 161558 76102
rect 161130 75922 161186 75978
rect 161254 75922 161310 75978
rect 161378 75922 161434 75978
rect 161502 75922 161558 75978
rect 161930 64294 161986 64350
rect 162054 64294 162110 64350
rect 162178 64294 162234 64350
rect 162302 64294 162358 64350
rect 161930 64170 161986 64226
rect 162054 64170 162110 64226
rect 162178 64170 162234 64226
rect 162302 64170 162358 64226
rect 161930 64046 161986 64102
rect 162054 64046 162110 64102
rect 162178 64046 162234 64102
rect 162302 64046 162358 64102
rect 161930 63922 161986 63978
rect 162054 63922 162110 63978
rect 162178 63922 162234 63978
rect 162302 63922 162358 63978
rect 162834 64294 162890 64350
rect 162958 64294 163014 64350
rect 163082 64294 163138 64350
rect 163206 64294 163262 64350
rect 162834 64170 162890 64226
rect 162958 64170 163014 64226
rect 163082 64170 163138 64226
rect 163206 64170 163262 64226
rect 162834 64046 162890 64102
rect 162958 64046 163014 64102
rect 163082 64046 163138 64102
rect 163206 64046 163262 64102
rect 162834 63922 162890 63978
rect 162958 63922 163014 63978
rect 163082 63922 163138 63978
rect 163206 63922 163262 63978
rect 161130 58294 161186 58350
rect 161254 58294 161310 58350
rect 161378 58294 161434 58350
rect 161502 58294 161558 58350
rect 161130 58170 161186 58226
rect 161254 58170 161310 58226
rect 161378 58170 161434 58226
rect 161502 58170 161558 58226
rect 161130 58046 161186 58102
rect 161254 58046 161310 58102
rect 161378 58046 161434 58102
rect 161502 58046 161558 58102
rect 161130 57922 161186 57978
rect 161254 57922 161310 57978
rect 161378 57922 161434 57978
rect 161502 57922 161558 57978
rect 161930 46294 161986 46350
rect 162054 46294 162110 46350
rect 162178 46294 162234 46350
rect 162302 46294 162358 46350
rect 161930 46170 161986 46226
rect 162054 46170 162110 46226
rect 162178 46170 162234 46226
rect 162302 46170 162358 46226
rect 161930 46046 161986 46102
rect 162054 46046 162110 46102
rect 162178 46046 162234 46102
rect 162302 46046 162358 46102
rect 161930 45922 161986 45978
rect 162054 45922 162110 45978
rect 162178 45922 162234 45978
rect 162302 45922 162358 45978
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 172038 190294 172094 190350
rect 172162 190294 172218 190350
rect 172038 190170 172094 190226
rect 172162 190170 172218 190226
rect 172038 190046 172094 190102
rect 172162 190046 172218 190102
rect 172038 189922 172094 189978
rect 172162 189922 172218 189978
rect 172038 172294 172094 172350
rect 172162 172294 172218 172350
rect 172038 172170 172094 172226
rect 172162 172170 172218 172226
rect 172038 172046 172094 172102
rect 172162 172046 172218 172102
rect 172038 171922 172094 171978
rect 172162 171922 172218 171978
rect 187398 202294 187454 202350
rect 187522 202294 187578 202350
rect 187398 202170 187454 202226
rect 187522 202170 187578 202226
rect 187398 202046 187454 202102
rect 187522 202046 187578 202102
rect 187398 201922 187454 201978
rect 187522 201922 187578 201978
rect 187398 184294 187454 184350
rect 187522 184294 187578 184350
rect 187398 184170 187454 184226
rect 187522 184170 187578 184226
rect 187398 184046 187454 184102
rect 187522 184046 187578 184102
rect 187398 183922 187454 183978
rect 187522 183922 187578 183978
rect 185612 175562 185668 175618
rect 187398 166294 187454 166350
rect 187522 166294 187578 166350
rect 187398 166170 187454 166226
rect 187522 166170 187578 166226
rect 187398 166046 187454 166102
rect 187522 166046 187578 166102
rect 187398 165922 187454 165978
rect 187522 165922 187578 165978
rect 193554 298294 193610 298350
rect 193678 298294 193734 298350
rect 193802 298294 193858 298350
rect 193926 298294 193982 298350
rect 193554 298170 193610 298226
rect 193678 298170 193734 298226
rect 193802 298170 193858 298226
rect 193926 298170 193982 298226
rect 193554 298046 193610 298102
rect 193678 298046 193734 298102
rect 193802 298046 193858 298102
rect 193926 298046 193982 298102
rect 193554 297922 193610 297978
rect 193678 297922 193734 297978
rect 193802 297922 193858 297978
rect 193926 297922 193982 297978
rect 189834 274294 189890 274350
rect 189958 274294 190014 274350
rect 190082 274294 190138 274350
rect 190206 274294 190262 274350
rect 189834 274170 189890 274226
rect 189958 274170 190014 274226
rect 190082 274170 190138 274226
rect 190206 274170 190262 274226
rect 189834 274046 189890 274102
rect 189958 274046 190014 274102
rect 190082 274046 190138 274102
rect 190206 274046 190262 274102
rect 189834 273922 189890 273978
rect 189958 273922 190014 273978
rect 190082 273922 190138 273978
rect 190206 273922 190262 273978
rect 189834 256294 189890 256350
rect 189958 256294 190014 256350
rect 190082 256294 190138 256350
rect 190206 256294 190262 256350
rect 189834 256170 189890 256226
rect 189958 256170 190014 256226
rect 190082 256170 190138 256226
rect 190206 256170 190262 256226
rect 189834 256046 189890 256102
rect 189958 256046 190014 256102
rect 190082 256046 190138 256102
rect 190206 256046 190262 256102
rect 189834 255922 189890 255978
rect 189958 255922 190014 255978
rect 190082 255922 190138 255978
rect 190206 255922 190262 255978
rect 189834 238294 189890 238350
rect 189958 238294 190014 238350
rect 190082 238294 190138 238350
rect 190206 238294 190262 238350
rect 189834 238170 189890 238226
rect 189958 238170 190014 238226
rect 190082 238170 190138 238226
rect 190206 238170 190262 238226
rect 189834 238046 189890 238102
rect 189958 238046 190014 238102
rect 190082 238046 190138 238102
rect 190206 238046 190262 238102
rect 189834 237922 189890 237978
rect 189958 237922 190014 237978
rect 190082 237922 190138 237978
rect 190206 237922 190262 237978
rect 189834 220294 189890 220350
rect 189958 220294 190014 220350
rect 190082 220294 190138 220350
rect 190206 220294 190262 220350
rect 189834 220170 189890 220226
rect 189958 220170 190014 220226
rect 190082 220170 190138 220226
rect 190206 220170 190262 220226
rect 189834 220046 189890 220102
rect 189958 220046 190014 220102
rect 190082 220046 190138 220102
rect 190206 220046 190262 220102
rect 189834 219922 189890 219978
rect 189958 219922 190014 219978
rect 190082 219922 190138 219978
rect 190206 219922 190262 219978
rect 189834 202294 189890 202350
rect 189958 202294 190014 202350
rect 190082 202294 190138 202350
rect 190206 202294 190262 202350
rect 189834 202170 189890 202226
rect 189958 202170 190014 202226
rect 190082 202170 190138 202226
rect 190206 202170 190262 202226
rect 189834 202046 189890 202102
rect 189958 202046 190014 202102
rect 190082 202046 190138 202102
rect 190206 202046 190262 202102
rect 189834 201922 189890 201978
rect 189958 201922 190014 201978
rect 190082 201922 190138 201978
rect 190206 201922 190262 201978
rect 189834 184294 189890 184350
rect 189958 184294 190014 184350
rect 190082 184294 190138 184350
rect 190206 184294 190262 184350
rect 189834 184170 189890 184226
rect 189958 184170 190014 184226
rect 190082 184170 190138 184226
rect 190206 184170 190262 184226
rect 189834 184046 189890 184102
rect 189958 184046 190014 184102
rect 190082 184046 190138 184102
rect 190206 184046 190262 184102
rect 189834 183922 189890 183978
rect 189958 183922 190014 183978
rect 190082 183922 190138 183978
rect 190206 183922 190262 183978
rect 188972 173942 189028 173998
rect 189834 166294 189890 166350
rect 189958 166294 190014 166350
rect 190082 166294 190138 166350
rect 190206 166294 190262 166350
rect 189834 166170 189890 166226
rect 189958 166170 190014 166226
rect 190082 166170 190138 166226
rect 190206 166170 190262 166226
rect 189834 166046 189890 166102
rect 189958 166046 190014 166102
rect 190082 166046 190138 166102
rect 190206 166046 190262 166102
rect 189834 165922 189890 165978
rect 189958 165922 190014 165978
rect 190082 165922 190138 165978
rect 190206 165922 190262 165978
rect 202758 298294 202814 298350
rect 202882 298294 202938 298350
rect 202758 298170 202814 298226
rect 202882 298170 202938 298226
rect 202758 298046 202814 298102
rect 202882 298046 202938 298102
rect 202758 297922 202814 297978
rect 202882 297922 202938 297978
rect 220554 292294 220610 292350
rect 220678 292294 220734 292350
rect 220802 292294 220858 292350
rect 220926 292294 220982 292350
rect 220554 292170 220610 292226
rect 220678 292170 220734 292226
rect 220802 292170 220858 292226
rect 220926 292170 220982 292226
rect 220554 292046 220610 292102
rect 220678 292046 220734 292102
rect 220802 292046 220858 292102
rect 220926 292046 220982 292102
rect 220554 291922 220610 291978
rect 220678 291922 220734 291978
rect 220802 291922 220858 291978
rect 220926 291922 220982 291978
rect 193554 280294 193610 280350
rect 193678 280294 193734 280350
rect 193802 280294 193858 280350
rect 193926 280294 193982 280350
rect 193554 280170 193610 280226
rect 193678 280170 193734 280226
rect 193802 280170 193858 280226
rect 193926 280170 193982 280226
rect 193554 280046 193610 280102
rect 193678 280046 193734 280102
rect 193802 280046 193858 280102
rect 193926 280046 193982 280102
rect 193554 279922 193610 279978
rect 193678 279922 193734 279978
rect 193802 279922 193858 279978
rect 193926 279922 193982 279978
rect 193554 262294 193610 262350
rect 193678 262294 193734 262350
rect 193802 262294 193858 262350
rect 193926 262294 193982 262350
rect 193554 262170 193610 262226
rect 193678 262170 193734 262226
rect 193802 262170 193858 262226
rect 193926 262170 193982 262226
rect 193554 262046 193610 262102
rect 193678 262046 193734 262102
rect 193802 262046 193858 262102
rect 193926 262046 193982 262102
rect 193554 261922 193610 261978
rect 193678 261922 193734 261978
rect 193802 261922 193858 261978
rect 193926 261922 193982 261978
rect 193554 244294 193610 244350
rect 193678 244294 193734 244350
rect 193802 244294 193858 244350
rect 193926 244294 193982 244350
rect 193554 244170 193610 244226
rect 193678 244170 193734 244226
rect 193802 244170 193858 244226
rect 193926 244170 193982 244226
rect 193554 244046 193610 244102
rect 193678 244046 193734 244102
rect 193802 244046 193858 244102
rect 193926 244046 193982 244102
rect 193554 243922 193610 243978
rect 193678 243922 193734 243978
rect 193802 243922 193858 243978
rect 193926 243922 193982 243978
rect 193554 226294 193610 226350
rect 193678 226294 193734 226350
rect 193802 226294 193858 226350
rect 193926 226294 193982 226350
rect 193554 226170 193610 226226
rect 193678 226170 193734 226226
rect 193802 226170 193858 226226
rect 193926 226170 193982 226226
rect 193554 226046 193610 226102
rect 193678 226046 193734 226102
rect 193802 226046 193858 226102
rect 193926 226046 193982 226102
rect 193554 225922 193610 225978
rect 193678 225922 193734 225978
rect 193802 225922 193858 225978
rect 193926 225922 193982 225978
rect 193554 208294 193610 208350
rect 193678 208294 193734 208350
rect 193802 208294 193858 208350
rect 193926 208294 193982 208350
rect 193554 208170 193610 208226
rect 193678 208170 193734 208226
rect 193802 208170 193858 208226
rect 193926 208170 193982 208226
rect 193554 208046 193610 208102
rect 193678 208046 193734 208102
rect 193802 208046 193858 208102
rect 193926 208046 193982 208102
rect 193554 207922 193610 207978
rect 193678 207922 193734 207978
rect 193802 207922 193858 207978
rect 193926 207922 193982 207978
rect 193554 190294 193610 190350
rect 193678 190294 193734 190350
rect 193802 190294 193858 190350
rect 193926 190294 193982 190350
rect 193554 190170 193610 190226
rect 193678 190170 193734 190226
rect 193802 190170 193858 190226
rect 193926 190170 193982 190226
rect 193554 190046 193610 190102
rect 193678 190046 193734 190102
rect 193802 190046 193858 190102
rect 193926 190046 193982 190102
rect 193554 189922 193610 189978
rect 193678 189922 193734 189978
rect 193802 189922 193858 189978
rect 193926 189922 193982 189978
rect 193554 172294 193610 172350
rect 193678 172294 193734 172350
rect 193802 172294 193858 172350
rect 193926 172294 193982 172350
rect 193554 172170 193610 172226
rect 193678 172170 193734 172226
rect 193802 172170 193858 172226
rect 193926 172170 193982 172226
rect 193554 172046 193610 172102
rect 193678 172046 193734 172102
rect 193802 172046 193858 172102
rect 193926 172046 193982 172102
rect 193554 171922 193610 171978
rect 193678 171922 193734 171978
rect 193802 171922 193858 171978
rect 193926 171922 193982 171978
rect 192332 170702 192388 170758
rect 189834 148294 189890 148350
rect 189958 148294 190014 148350
rect 190082 148294 190138 148350
rect 190206 148294 190262 148350
rect 189834 148170 189890 148226
rect 189958 148170 190014 148226
rect 190082 148170 190138 148226
rect 190206 148170 190262 148226
rect 189834 148046 189890 148102
rect 189958 148046 190014 148102
rect 190082 148046 190138 148102
rect 190206 148046 190262 148102
rect 189834 147922 189890 147978
rect 189958 147922 190014 147978
rect 190082 147922 190138 147978
rect 190206 147922 190262 147978
rect 189834 130294 189890 130350
rect 189958 130294 190014 130350
rect 190082 130294 190138 130350
rect 190206 130294 190262 130350
rect 189834 130170 189890 130226
rect 189958 130170 190014 130226
rect 190082 130170 190138 130226
rect 190206 130170 190262 130226
rect 189834 130046 189890 130102
rect 189958 130046 190014 130102
rect 190082 130046 190138 130102
rect 190206 130046 190262 130102
rect 189834 129922 189890 129978
rect 189958 129922 190014 129978
rect 190082 129922 190138 129978
rect 190206 129922 190262 129978
rect 189834 112294 189890 112350
rect 189958 112294 190014 112350
rect 190082 112294 190138 112350
rect 190206 112294 190262 112350
rect 189834 112170 189890 112226
rect 189958 112170 190014 112226
rect 190082 112170 190138 112226
rect 190206 112170 190262 112226
rect 189834 112046 189890 112102
rect 189958 112046 190014 112102
rect 190082 112046 190138 112102
rect 190206 112046 190262 112102
rect 189834 111922 189890 111978
rect 189958 111922 190014 111978
rect 190082 111922 190138 111978
rect 190206 111922 190262 111978
rect 189834 94294 189890 94350
rect 189958 94294 190014 94350
rect 190082 94294 190138 94350
rect 190206 94294 190262 94350
rect 189834 94170 189890 94226
rect 189958 94170 190014 94226
rect 190082 94170 190138 94226
rect 190206 94170 190262 94226
rect 189834 94046 189890 94102
rect 189958 94046 190014 94102
rect 190082 94046 190138 94102
rect 190206 94046 190262 94102
rect 189834 93922 189890 93978
rect 189958 93922 190014 93978
rect 190082 93922 190138 93978
rect 190206 93922 190262 93978
rect 189834 76294 189890 76350
rect 189958 76294 190014 76350
rect 190082 76294 190138 76350
rect 190206 76294 190262 76350
rect 189834 76170 189890 76226
rect 189958 76170 190014 76226
rect 190082 76170 190138 76226
rect 190206 76170 190262 76226
rect 189834 76046 189890 76102
rect 189958 76046 190014 76102
rect 190082 76046 190138 76102
rect 190206 76046 190262 76102
rect 189834 75922 189890 75978
rect 189958 75922 190014 75978
rect 190082 75922 190138 75978
rect 190206 75922 190262 75978
rect 189834 58294 189890 58350
rect 189958 58294 190014 58350
rect 190082 58294 190138 58350
rect 190206 58294 190262 58350
rect 189834 58170 189890 58226
rect 189958 58170 190014 58226
rect 190082 58170 190138 58226
rect 190206 58170 190262 58226
rect 189834 58046 189890 58102
rect 189958 58046 190014 58102
rect 190082 58046 190138 58102
rect 190206 58046 190262 58102
rect 189834 57922 189890 57978
rect 189958 57922 190014 57978
rect 190082 57922 190138 57978
rect 190206 57922 190262 57978
rect 189834 40294 189890 40350
rect 189958 40294 190014 40350
rect 190082 40294 190138 40350
rect 190206 40294 190262 40350
rect 189834 40170 189890 40226
rect 189958 40170 190014 40226
rect 190082 40170 190138 40226
rect 190206 40170 190262 40226
rect 189834 40046 189890 40102
rect 189958 40046 190014 40102
rect 190082 40046 190138 40102
rect 190206 40046 190262 40102
rect 189834 39922 189890 39978
rect 189958 39922 190014 39978
rect 190082 39922 190138 39978
rect 190206 39922 190262 39978
rect 189834 22294 189890 22350
rect 189958 22294 190014 22350
rect 190082 22294 190138 22350
rect 190206 22294 190262 22350
rect 189834 22170 189890 22226
rect 189958 22170 190014 22226
rect 190082 22170 190138 22226
rect 190206 22170 190262 22226
rect 189834 22046 189890 22102
rect 189958 22046 190014 22102
rect 190082 22046 190138 22102
rect 190206 22046 190262 22102
rect 189834 21922 189890 21978
rect 189958 21922 190014 21978
rect 190082 21922 190138 21978
rect 190206 21922 190262 21978
rect 193554 154294 193610 154350
rect 193678 154294 193734 154350
rect 193802 154294 193858 154350
rect 193926 154294 193982 154350
rect 193554 154170 193610 154226
rect 193678 154170 193734 154226
rect 193802 154170 193858 154226
rect 193926 154170 193982 154226
rect 193554 154046 193610 154102
rect 193678 154046 193734 154102
rect 193802 154046 193858 154102
rect 193926 154046 193982 154102
rect 193554 153922 193610 153978
rect 193678 153922 193734 153978
rect 193802 153922 193858 153978
rect 193926 153922 193982 153978
rect 195692 168902 195748 168958
rect 193554 136294 193610 136350
rect 193678 136294 193734 136350
rect 193802 136294 193858 136350
rect 193926 136294 193982 136350
rect 193554 136170 193610 136226
rect 193678 136170 193734 136226
rect 193802 136170 193858 136226
rect 193926 136170 193982 136226
rect 193554 136046 193610 136102
rect 193678 136046 193734 136102
rect 193802 136046 193858 136102
rect 193926 136046 193982 136102
rect 193554 135922 193610 135978
rect 193678 135922 193734 135978
rect 193802 135922 193858 135978
rect 193926 135922 193982 135978
rect 193554 118294 193610 118350
rect 193678 118294 193734 118350
rect 193802 118294 193858 118350
rect 193926 118294 193982 118350
rect 193554 118170 193610 118226
rect 193678 118170 193734 118226
rect 193802 118170 193858 118226
rect 193926 118170 193982 118226
rect 193554 118046 193610 118102
rect 193678 118046 193734 118102
rect 193802 118046 193858 118102
rect 193926 118046 193982 118102
rect 193554 117922 193610 117978
rect 193678 117922 193734 117978
rect 193802 117922 193858 117978
rect 193926 117922 193982 117978
rect 193554 100294 193610 100350
rect 193678 100294 193734 100350
rect 193802 100294 193858 100350
rect 193926 100294 193982 100350
rect 193554 100170 193610 100226
rect 193678 100170 193734 100226
rect 193802 100170 193858 100226
rect 193926 100170 193982 100226
rect 193554 100046 193610 100102
rect 193678 100046 193734 100102
rect 193802 100046 193858 100102
rect 193926 100046 193982 100102
rect 193554 99922 193610 99978
rect 193678 99922 193734 99978
rect 193802 99922 193858 99978
rect 193926 99922 193982 99978
rect 193554 82294 193610 82350
rect 193678 82294 193734 82350
rect 193802 82294 193858 82350
rect 193926 82294 193982 82350
rect 193554 82170 193610 82226
rect 193678 82170 193734 82226
rect 193802 82170 193858 82226
rect 193926 82170 193982 82226
rect 193554 82046 193610 82102
rect 193678 82046 193734 82102
rect 193802 82046 193858 82102
rect 193926 82046 193982 82102
rect 193554 81922 193610 81978
rect 193678 81922 193734 81978
rect 193802 81922 193858 81978
rect 193926 81922 193982 81978
rect 193554 64294 193610 64350
rect 193678 64294 193734 64350
rect 193802 64294 193858 64350
rect 193926 64294 193982 64350
rect 193554 64170 193610 64226
rect 193678 64170 193734 64226
rect 193802 64170 193858 64226
rect 193926 64170 193982 64226
rect 193554 64046 193610 64102
rect 193678 64046 193734 64102
rect 193802 64046 193858 64102
rect 193926 64046 193982 64102
rect 193554 63922 193610 63978
rect 193678 63922 193734 63978
rect 193802 63922 193858 63978
rect 193926 63922 193982 63978
rect 193554 46294 193610 46350
rect 193678 46294 193734 46350
rect 193802 46294 193858 46350
rect 193926 46294 193982 46350
rect 193554 46170 193610 46226
rect 193678 46170 193734 46226
rect 193802 46170 193858 46226
rect 193926 46170 193982 46226
rect 193554 46046 193610 46102
rect 193678 46046 193734 46102
rect 193802 46046 193858 46102
rect 193926 46046 193982 46102
rect 193554 45922 193610 45978
rect 193678 45922 193734 45978
rect 193802 45922 193858 45978
rect 193926 45922 193982 45978
rect 193554 28294 193610 28350
rect 193678 28294 193734 28350
rect 193802 28294 193858 28350
rect 193926 28294 193982 28350
rect 193554 28170 193610 28226
rect 193678 28170 193734 28226
rect 193802 28170 193858 28226
rect 193926 28170 193982 28226
rect 193554 28046 193610 28102
rect 193678 28046 193734 28102
rect 193802 28046 193858 28102
rect 193926 28046 193982 28102
rect 193554 27922 193610 27978
rect 193678 27922 193734 27978
rect 193802 27922 193858 27978
rect 193926 27922 193982 27978
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 202758 190294 202814 190350
rect 202882 190294 202938 190350
rect 202758 190170 202814 190226
rect 202882 190170 202938 190226
rect 202758 190046 202814 190102
rect 202882 190046 202938 190102
rect 202758 189922 202814 189978
rect 202882 189922 202938 189978
rect 203308 173762 203364 173818
rect 202758 172294 202814 172350
rect 202882 172294 202938 172350
rect 202758 172170 202814 172226
rect 202882 172170 202938 172226
rect 202758 172046 202814 172102
rect 202882 172046 202938 172102
rect 202758 171922 202814 171978
rect 202882 171922 202938 171978
rect 200732 170522 200788 170578
rect 218118 202294 218174 202350
rect 218242 202294 218298 202350
rect 218118 202170 218174 202226
rect 218242 202170 218298 202226
rect 218118 202046 218174 202102
rect 218242 202046 218298 202102
rect 218118 201922 218174 201978
rect 218242 201922 218298 201978
rect 218118 184294 218174 184350
rect 218242 184294 218298 184350
rect 218118 184170 218174 184226
rect 218242 184170 218298 184226
rect 218118 184046 218174 184102
rect 218242 184046 218298 184102
rect 218118 183922 218174 183978
rect 218242 183922 218298 183978
rect 218428 175562 218484 175618
rect 224274 298294 224330 298350
rect 224398 298294 224454 298350
rect 224522 298294 224578 298350
rect 224646 298294 224702 298350
rect 224274 298170 224330 298226
rect 224398 298170 224454 298226
rect 224522 298170 224578 298226
rect 224646 298170 224702 298226
rect 224274 298046 224330 298102
rect 224398 298046 224454 298102
rect 224522 298046 224578 298102
rect 224646 298046 224702 298102
rect 224274 297922 224330 297978
rect 224398 297922 224454 297978
rect 224522 297922 224578 297978
rect 224646 297922 224702 297978
rect 220554 274294 220610 274350
rect 220678 274294 220734 274350
rect 220802 274294 220858 274350
rect 220926 274294 220982 274350
rect 220554 274170 220610 274226
rect 220678 274170 220734 274226
rect 220802 274170 220858 274226
rect 220926 274170 220982 274226
rect 220554 274046 220610 274102
rect 220678 274046 220734 274102
rect 220802 274046 220858 274102
rect 220926 274046 220982 274102
rect 220554 273922 220610 273978
rect 220678 273922 220734 273978
rect 220802 273922 220858 273978
rect 220926 273922 220982 273978
rect 220554 256294 220610 256350
rect 220678 256294 220734 256350
rect 220802 256294 220858 256350
rect 220926 256294 220982 256350
rect 220554 256170 220610 256226
rect 220678 256170 220734 256226
rect 220802 256170 220858 256226
rect 220926 256170 220982 256226
rect 220554 256046 220610 256102
rect 220678 256046 220734 256102
rect 220802 256046 220858 256102
rect 220926 256046 220982 256102
rect 220554 255922 220610 255978
rect 220678 255922 220734 255978
rect 220802 255922 220858 255978
rect 220926 255922 220982 255978
rect 220554 238294 220610 238350
rect 220678 238294 220734 238350
rect 220802 238294 220858 238350
rect 220926 238294 220982 238350
rect 220554 238170 220610 238226
rect 220678 238170 220734 238226
rect 220802 238170 220858 238226
rect 220926 238170 220982 238226
rect 220554 238046 220610 238102
rect 220678 238046 220734 238102
rect 220802 238046 220858 238102
rect 220926 238046 220982 238102
rect 220554 237922 220610 237978
rect 220678 237922 220734 237978
rect 220802 237922 220858 237978
rect 220926 237922 220982 237978
rect 220554 220294 220610 220350
rect 220678 220294 220734 220350
rect 220802 220294 220858 220350
rect 220926 220294 220982 220350
rect 220554 220170 220610 220226
rect 220678 220170 220734 220226
rect 220802 220170 220858 220226
rect 220926 220170 220982 220226
rect 220554 220046 220610 220102
rect 220678 220046 220734 220102
rect 220802 220046 220858 220102
rect 220926 220046 220982 220102
rect 220554 219922 220610 219978
rect 220678 219922 220734 219978
rect 220802 219922 220858 219978
rect 220926 219922 220982 219978
rect 220554 202294 220610 202350
rect 220678 202294 220734 202350
rect 220802 202294 220858 202350
rect 220926 202294 220982 202350
rect 220554 202170 220610 202226
rect 220678 202170 220734 202226
rect 220802 202170 220858 202226
rect 220926 202170 220982 202226
rect 220554 202046 220610 202102
rect 220678 202046 220734 202102
rect 220802 202046 220858 202102
rect 220926 202046 220982 202102
rect 220554 201922 220610 201978
rect 220678 201922 220734 201978
rect 220802 201922 220858 201978
rect 220926 201922 220982 201978
rect 220554 184294 220610 184350
rect 220678 184294 220734 184350
rect 220802 184294 220858 184350
rect 220926 184294 220982 184350
rect 220554 184170 220610 184226
rect 220678 184170 220734 184226
rect 220802 184170 220858 184226
rect 220926 184170 220982 184226
rect 220554 184046 220610 184102
rect 220678 184046 220734 184102
rect 220802 184046 220858 184102
rect 220926 184046 220982 184102
rect 220554 183922 220610 183978
rect 220678 183922 220734 183978
rect 220802 183922 220858 183978
rect 220926 183922 220982 183978
rect 215068 170702 215124 170758
rect 221788 173942 221844 173998
rect 233478 298294 233534 298350
rect 233602 298294 233658 298350
rect 233478 298170 233534 298226
rect 233602 298170 233658 298226
rect 233478 298046 233534 298102
rect 233602 298046 233658 298102
rect 233478 297922 233534 297978
rect 233602 297922 233658 297978
rect 251274 292294 251330 292350
rect 251398 292294 251454 292350
rect 251522 292294 251578 292350
rect 251646 292294 251702 292350
rect 251274 292170 251330 292226
rect 251398 292170 251454 292226
rect 251522 292170 251578 292226
rect 251646 292170 251702 292226
rect 251274 292046 251330 292102
rect 251398 292046 251454 292102
rect 251522 292046 251578 292102
rect 251646 292046 251702 292102
rect 251274 291922 251330 291978
rect 251398 291922 251454 291978
rect 251522 291922 251578 291978
rect 251646 291922 251702 291978
rect 224274 280294 224330 280350
rect 224398 280294 224454 280350
rect 224522 280294 224578 280350
rect 224646 280294 224702 280350
rect 224274 280170 224330 280226
rect 224398 280170 224454 280226
rect 224522 280170 224578 280226
rect 224646 280170 224702 280226
rect 224274 280046 224330 280102
rect 224398 280046 224454 280102
rect 224522 280046 224578 280102
rect 224646 280046 224702 280102
rect 224274 279922 224330 279978
rect 224398 279922 224454 279978
rect 224522 279922 224578 279978
rect 224646 279922 224702 279978
rect 224274 262294 224330 262350
rect 224398 262294 224454 262350
rect 224522 262294 224578 262350
rect 224646 262294 224702 262350
rect 224274 262170 224330 262226
rect 224398 262170 224454 262226
rect 224522 262170 224578 262226
rect 224646 262170 224702 262226
rect 224274 262046 224330 262102
rect 224398 262046 224454 262102
rect 224522 262046 224578 262102
rect 224646 262046 224702 262102
rect 224274 261922 224330 261978
rect 224398 261922 224454 261978
rect 224522 261922 224578 261978
rect 224646 261922 224702 261978
rect 224274 244294 224330 244350
rect 224398 244294 224454 244350
rect 224522 244294 224578 244350
rect 224646 244294 224702 244350
rect 224274 244170 224330 244226
rect 224398 244170 224454 244226
rect 224522 244170 224578 244226
rect 224646 244170 224702 244226
rect 224274 244046 224330 244102
rect 224398 244046 224454 244102
rect 224522 244046 224578 244102
rect 224646 244046 224702 244102
rect 224274 243922 224330 243978
rect 224398 243922 224454 243978
rect 224522 243922 224578 243978
rect 224646 243922 224702 243978
rect 224274 226294 224330 226350
rect 224398 226294 224454 226350
rect 224522 226294 224578 226350
rect 224646 226294 224702 226350
rect 224274 226170 224330 226226
rect 224398 226170 224454 226226
rect 224522 226170 224578 226226
rect 224646 226170 224702 226226
rect 224274 226046 224330 226102
rect 224398 226046 224454 226102
rect 224522 226046 224578 226102
rect 224646 226046 224702 226102
rect 224274 225922 224330 225978
rect 224398 225922 224454 225978
rect 224522 225922 224578 225978
rect 224646 225922 224702 225978
rect 224274 208294 224330 208350
rect 224398 208294 224454 208350
rect 224522 208294 224578 208350
rect 224646 208294 224702 208350
rect 224274 208170 224330 208226
rect 224398 208170 224454 208226
rect 224522 208170 224578 208226
rect 224646 208170 224702 208226
rect 224274 208046 224330 208102
rect 224398 208046 224454 208102
rect 224522 208046 224578 208102
rect 224646 208046 224702 208102
rect 224274 207922 224330 207978
rect 224398 207922 224454 207978
rect 224522 207922 224578 207978
rect 224646 207922 224702 207978
rect 224274 190294 224330 190350
rect 224398 190294 224454 190350
rect 224522 190294 224578 190350
rect 224646 190294 224702 190350
rect 224274 190170 224330 190226
rect 224398 190170 224454 190226
rect 224522 190170 224578 190226
rect 224646 190170 224702 190226
rect 224274 190046 224330 190102
rect 224398 190046 224454 190102
rect 224522 190046 224578 190102
rect 224646 190046 224702 190102
rect 224274 189922 224330 189978
rect 224398 189922 224454 189978
rect 224522 189922 224578 189978
rect 224646 189922 224702 189978
rect 224274 172294 224330 172350
rect 224398 172294 224454 172350
rect 224522 172294 224578 172350
rect 224646 172294 224702 172350
rect 224274 172170 224330 172226
rect 224398 172170 224454 172226
rect 224522 172170 224578 172226
rect 224646 172170 224702 172226
rect 224274 172046 224330 172102
rect 224398 172046 224454 172102
rect 224522 172046 224578 172102
rect 224646 172046 224702 172102
rect 224274 171922 224330 171978
rect 224398 171922 224454 171978
rect 224522 171922 224578 171978
rect 224646 171922 224702 171978
rect 213388 168902 213444 168958
rect 208348 168722 208404 168778
rect 198268 167282 198324 167338
rect 218118 166294 218174 166350
rect 218242 166294 218298 166350
rect 218118 166170 218174 166226
rect 218242 166170 218298 166226
rect 218118 166046 218174 166102
rect 218242 166046 218298 166102
rect 218118 165922 218174 165978
rect 218242 165922 218298 165978
rect 220554 148294 220610 148350
rect 220678 148294 220734 148350
rect 220802 148294 220858 148350
rect 220926 148294 220982 148350
rect 220554 148170 220610 148226
rect 220678 148170 220734 148226
rect 220802 148170 220858 148226
rect 220926 148170 220982 148226
rect 220554 148046 220610 148102
rect 220678 148046 220734 148102
rect 220802 148046 220858 148102
rect 220926 148046 220982 148102
rect 220554 147922 220610 147978
rect 220678 147922 220734 147978
rect 220802 147922 220858 147978
rect 220926 147922 220982 147978
rect 219324 141902 219380 141958
rect 214620 141002 214676 141058
rect 220554 130294 220610 130350
rect 220678 130294 220734 130350
rect 220802 130294 220858 130350
rect 220926 130294 220982 130350
rect 220554 130170 220610 130226
rect 220678 130170 220734 130226
rect 220802 130170 220858 130226
rect 220926 130170 220982 130226
rect 220554 130046 220610 130102
rect 220678 130046 220734 130102
rect 220802 130046 220858 130102
rect 220926 130046 220982 130102
rect 220554 129922 220610 129978
rect 220678 129922 220734 129978
rect 220802 129922 220858 129978
rect 220926 129922 220982 129978
rect 220554 112294 220610 112350
rect 220678 112294 220734 112350
rect 220802 112294 220858 112350
rect 220926 112294 220982 112350
rect 220554 112170 220610 112226
rect 220678 112170 220734 112226
rect 220802 112170 220858 112226
rect 220926 112170 220982 112226
rect 220554 112046 220610 112102
rect 220678 112046 220734 112102
rect 220802 112046 220858 112102
rect 220926 112046 220982 112102
rect 220554 111922 220610 111978
rect 220678 111922 220734 111978
rect 220802 111922 220858 111978
rect 220926 111922 220982 111978
rect 220554 94294 220610 94350
rect 220678 94294 220734 94350
rect 220802 94294 220858 94350
rect 220926 94294 220982 94350
rect 220554 94170 220610 94226
rect 220678 94170 220734 94226
rect 220802 94170 220858 94226
rect 220926 94170 220982 94226
rect 220554 94046 220610 94102
rect 220678 94046 220734 94102
rect 220802 94046 220858 94102
rect 220926 94046 220982 94102
rect 220554 93922 220610 93978
rect 220678 93922 220734 93978
rect 220802 93922 220858 93978
rect 220926 93922 220982 93978
rect 220554 76294 220610 76350
rect 220678 76294 220734 76350
rect 220802 76294 220858 76350
rect 220926 76294 220982 76350
rect 220554 76170 220610 76226
rect 220678 76170 220734 76226
rect 220802 76170 220858 76226
rect 220926 76170 220982 76226
rect 220554 76046 220610 76102
rect 220678 76046 220734 76102
rect 220802 76046 220858 76102
rect 220926 76046 220982 76102
rect 220554 75922 220610 75978
rect 220678 75922 220734 75978
rect 220802 75922 220858 75978
rect 220926 75922 220982 75978
rect 220554 58294 220610 58350
rect 220678 58294 220734 58350
rect 220802 58294 220858 58350
rect 220926 58294 220982 58350
rect 220554 58170 220610 58226
rect 220678 58170 220734 58226
rect 220802 58170 220858 58226
rect 220926 58170 220982 58226
rect 220554 58046 220610 58102
rect 220678 58046 220734 58102
rect 220802 58046 220858 58102
rect 220926 58046 220982 58102
rect 220554 57922 220610 57978
rect 220678 57922 220734 57978
rect 220802 57922 220858 57978
rect 220926 57922 220982 57978
rect 220554 40294 220610 40350
rect 220678 40294 220734 40350
rect 220802 40294 220858 40350
rect 220926 40294 220982 40350
rect 220554 40170 220610 40226
rect 220678 40170 220734 40226
rect 220802 40170 220858 40226
rect 220926 40170 220982 40226
rect 220554 40046 220610 40102
rect 220678 40046 220734 40102
rect 220802 40046 220858 40102
rect 220926 40046 220982 40102
rect 220554 39922 220610 39978
rect 220678 39922 220734 39978
rect 220802 39922 220858 39978
rect 220926 39922 220982 39978
rect 220554 22294 220610 22350
rect 220678 22294 220734 22350
rect 220802 22294 220858 22350
rect 220926 22294 220982 22350
rect 220554 22170 220610 22226
rect 220678 22170 220734 22226
rect 220802 22170 220858 22226
rect 220926 22170 220982 22226
rect 220554 22046 220610 22102
rect 220678 22046 220734 22102
rect 220802 22046 220858 22102
rect 220926 22046 220982 22102
rect 220554 21922 220610 21978
rect 220678 21922 220734 21978
rect 220802 21922 220858 21978
rect 220926 21922 220982 21978
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 224274 154294 224330 154350
rect 224398 154294 224454 154350
rect 224522 154294 224578 154350
rect 224646 154294 224702 154350
rect 224274 154170 224330 154226
rect 224398 154170 224454 154226
rect 224522 154170 224578 154226
rect 224646 154170 224702 154226
rect 224274 154046 224330 154102
rect 224398 154046 224454 154102
rect 224522 154046 224578 154102
rect 224646 154046 224702 154102
rect 224274 153922 224330 153978
rect 224398 153922 224454 153978
rect 224522 153922 224578 153978
rect 224646 153922 224702 153978
rect 224274 136294 224330 136350
rect 224398 136294 224454 136350
rect 224522 136294 224578 136350
rect 224646 136294 224702 136350
rect 224274 136170 224330 136226
rect 224398 136170 224454 136226
rect 224522 136170 224578 136226
rect 224646 136170 224702 136226
rect 224274 136046 224330 136102
rect 224398 136046 224454 136102
rect 224522 136046 224578 136102
rect 224646 136046 224702 136102
rect 224274 135922 224330 135978
rect 224398 135922 224454 135978
rect 224522 135922 224578 135978
rect 224646 135922 224702 135978
rect 224274 118294 224330 118350
rect 224398 118294 224454 118350
rect 224522 118294 224578 118350
rect 224646 118294 224702 118350
rect 224274 118170 224330 118226
rect 224398 118170 224454 118226
rect 224522 118170 224578 118226
rect 224646 118170 224702 118226
rect 224274 118046 224330 118102
rect 224398 118046 224454 118102
rect 224522 118046 224578 118102
rect 224646 118046 224702 118102
rect 224274 117922 224330 117978
rect 224398 117922 224454 117978
rect 224522 117922 224578 117978
rect 224646 117922 224702 117978
rect 224274 100294 224330 100350
rect 224398 100294 224454 100350
rect 224522 100294 224578 100350
rect 224646 100294 224702 100350
rect 224274 100170 224330 100226
rect 224398 100170 224454 100226
rect 224522 100170 224578 100226
rect 224646 100170 224702 100226
rect 224274 100046 224330 100102
rect 224398 100046 224454 100102
rect 224522 100046 224578 100102
rect 224646 100046 224702 100102
rect 224274 99922 224330 99978
rect 224398 99922 224454 99978
rect 224522 99922 224578 99978
rect 224646 99922 224702 99978
rect 224274 82294 224330 82350
rect 224398 82294 224454 82350
rect 224522 82294 224578 82350
rect 224646 82294 224702 82350
rect 224274 82170 224330 82226
rect 224398 82170 224454 82226
rect 224522 82170 224578 82226
rect 224646 82170 224702 82226
rect 224274 82046 224330 82102
rect 224398 82046 224454 82102
rect 224522 82046 224578 82102
rect 224646 82046 224702 82102
rect 224274 81922 224330 81978
rect 224398 81922 224454 81978
rect 224522 81922 224578 81978
rect 224646 81922 224702 81978
rect 224274 64294 224330 64350
rect 224398 64294 224454 64350
rect 224522 64294 224578 64350
rect 224646 64294 224702 64350
rect 224274 64170 224330 64226
rect 224398 64170 224454 64226
rect 224522 64170 224578 64226
rect 224646 64170 224702 64226
rect 224274 64046 224330 64102
rect 224398 64046 224454 64102
rect 224522 64046 224578 64102
rect 224646 64046 224702 64102
rect 224274 63922 224330 63978
rect 224398 63922 224454 63978
rect 224522 63922 224578 63978
rect 224646 63922 224702 63978
rect 224274 46294 224330 46350
rect 224398 46294 224454 46350
rect 224522 46294 224578 46350
rect 224646 46294 224702 46350
rect 224274 46170 224330 46226
rect 224398 46170 224454 46226
rect 224522 46170 224578 46226
rect 224646 46170 224702 46226
rect 224274 46046 224330 46102
rect 224398 46046 224454 46102
rect 224522 46046 224578 46102
rect 224646 46046 224702 46102
rect 224274 45922 224330 45978
rect 224398 45922 224454 45978
rect 224522 45922 224578 45978
rect 224646 45922 224702 45978
rect 224274 28294 224330 28350
rect 224398 28294 224454 28350
rect 224522 28294 224578 28350
rect 224646 28294 224702 28350
rect 224274 28170 224330 28226
rect 224398 28170 224454 28226
rect 224522 28170 224578 28226
rect 224646 28170 224702 28226
rect 224274 28046 224330 28102
rect 224398 28046 224454 28102
rect 224522 28046 224578 28102
rect 224646 28046 224702 28102
rect 224274 27922 224330 27978
rect 224398 27922 224454 27978
rect 224522 27922 224578 27978
rect 224646 27922 224702 27978
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 233478 190294 233534 190350
rect 233602 190294 233658 190350
rect 233478 190170 233534 190226
rect 233602 190170 233658 190226
rect 233478 190046 233534 190102
rect 233602 190046 233658 190102
rect 233478 189922 233534 189978
rect 233602 189922 233658 189978
rect 233478 172294 233534 172350
rect 233602 172294 233658 172350
rect 233478 172170 233534 172226
rect 233602 172170 233658 172226
rect 233478 172046 233534 172102
rect 233602 172046 233658 172102
rect 233478 171922 233534 171978
rect 233602 171922 233658 171978
rect 244636 142082 244692 142138
rect 245420 140822 245476 140878
rect 245812 130294 245868 130350
rect 245936 130294 245992 130350
rect 246060 130294 246116 130350
rect 246184 130294 246240 130350
rect 245812 130170 245868 130226
rect 245936 130170 245992 130226
rect 246060 130170 246116 130226
rect 246184 130170 246240 130226
rect 245812 130046 245868 130102
rect 245936 130046 245992 130102
rect 246060 130046 246116 130102
rect 246184 130046 246240 130102
rect 245812 129922 245868 129978
rect 245936 129922 245992 129978
rect 246060 129922 246116 129978
rect 246184 129922 246240 129978
rect 246612 118294 246668 118350
rect 246736 118294 246792 118350
rect 246860 118294 246916 118350
rect 246984 118294 247040 118350
rect 246612 118170 246668 118226
rect 246736 118170 246792 118226
rect 246860 118170 246916 118226
rect 246984 118170 247040 118226
rect 246612 118046 246668 118102
rect 246736 118046 246792 118102
rect 246860 118046 246916 118102
rect 246984 118046 247040 118102
rect 246612 117922 246668 117978
rect 246736 117922 246792 117978
rect 246860 117922 246916 117978
rect 246984 117922 247040 117978
rect 245812 112294 245868 112350
rect 245936 112294 245992 112350
rect 246060 112294 246116 112350
rect 246184 112294 246240 112350
rect 245812 112170 245868 112226
rect 245936 112170 245992 112226
rect 246060 112170 246116 112226
rect 246184 112170 246240 112226
rect 245812 112046 245868 112102
rect 245936 112046 245992 112102
rect 246060 112046 246116 112102
rect 246184 112046 246240 112102
rect 245812 111922 245868 111978
rect 245936 111922 245992 111978
rect 246060 111922 246116 111978
rect 246184 111922 246240 111978
rect 246612 100294 246668 100350
rect 246736 100294 246792 100350
rect 246860 100294 246916 100350
rect 246984 100294 247040 100350
rect 246612 100170 246668 100226
rect 246736 100170 246792 100226
rect 246860 100170 246916 100226
rect 246984 100170 247040 100226
rect 246612 100046 246668 100102
rect 246736 100046 246792 100102
rect 246860 100046 246916 100102
rect 246984 100046 247040 100102
rect 246612 99922 246668 99978
rect 246736 99922 246792 99978
rect 246860 99922 246916 99978
rect 246984 99922 247040 99978
rect 245812 94294 245868 94350
rect 245936 94294 245992 94350
rect 246060 94294 246116 94350
rect 246184 94294 246240 94350
rect 245812 94170 245868 94226
rect 245936 94170 245992 94226
rect 246060 94170 246116 94226
rect 246184 94170 246240 94226
rect 245812 94046 245868 94102
rect 245936 94046 245992 94102
rect 246060 94046 246116 94102
rect 246184 94046 246240 94102
rect 245812 93922 245868 93978
rect 245936 93922 245992 93978
rect 246060 93922 246116 93978
rect 246184 93922 246240 93978
rect 246612 82294 246668 82350
rect 246736 82294 246792 82350
rect 246860 82294 246916 82350
rect 246984 82294 247040 82350
rect 246612 82170 246668 82226
rect 246736 82170 246792 82226
rect 246860 82170 246916 82226
rect 246984 82170 247040 82226
rect 246612 82046 246668 82102
rect 246736 82046 246792 82102
rect 246860 82046 246916 82102
rect 246984 82046 247040 82102
rect 246612 81922 246668 81978
rect 246736 81922 246792 81978
rect 246860 81922 246916 81978
rect 246984 81922 247040 81978
rect 245812 76294 245868 76350
rect 245936 76294 245992 76350
rect 246060 76294 246116 76350
rect 246184 76294 246240 76350
rect 245812 76170 245868 76226
rect 245936 76170 245992 76226
rect 246060 76170 246116 76226
rect 246184 76170 246240 76226
rect 245812 76046 245868 76102
rect 245936 76046 245992 76102
rect 246060 76046 246116 76102
rect 246184 76046 246240 76102
rect 245812 75922 245868 75978
rect 245936 75922 245992 75978
rect 246060 75922 246116 75978
rect 246184 75922 246240 75978
rect 246612 64294 246668 64350
rect 246736 64294 246792 64350
rect 246860 64294 246916 64350
rect 246984 64294 247040 64350
rect 246612 64170 246668 64226
rect 246736 64170 246792 64226
rect 246860 64170 246916 64226
rect 246984 64170 247040 64226
rect 246612 64046 246668 64102
rect 246736 64046 246792 64102
rect 246860 64046 246916 64102
rect 246984 64046 247040 64102
rect 246612 63922 246668 63978
rect 246736 63922 246792 63978
rect 246860 63922 246916 63978
rect 246984 63922 247040 63978
rect 245812 58294 245868 58350
rect 245936 58294 245992 58350
rect 246060 58294 246116 58350
rect 246184 58294 246240 58350
rect 245812 58170 245868 58226
rect 245936 58170 245992 58226
rect 246060 58170 246116 58226
rect 246184 58170 246240 58226
rect 245812 58046 245868 58102
rect 245936 58046 245992 58102
rect 246060 58046 246116 58102
rect 246184 58046 246240 58102
rect 245812 57922 245868 57978
rect 245936 57922 245992 57978
rect 246060 57922 246116 57978
rect 246184 57922 246240 57978
rect 246612 46294 246668 46350
rect 246736 46294 246792 46350
rect 246860 46294 246916 46350
rect 246984 46294 247040 46350
rect 246612 46170 246668 46226
rect 246736 46170 246792 46226
rect 246860 46170 246916 46226
rect 246984 46170 247040 46226
rect 246612 46046 246668 46102
rect 246736 46046 246792 46102
rect 246860 46046 246916 46102
rect 246984 46046 247040 46102
rect 246612 45922 246668 45978
rect 246736 45922 246792 45978
rect 246860 45922 246916 45978
rect 246984 45922 247040 45978
rect 248838 202294 248894 202350
rect 248962 202294 249018 202350
rect 248838 202170 248894 202226
rect 248962 202170 249018 202226
rect 248838 202046 248894 202102
rect 248962 202046 249018 202102
rect 248838 201922 248894 201978
rect 248962 201922 249018 201978
rect 248838 184294 248894 184350
rect 248962 184294 249018 184350
rect 248838 184170 248894 184226
rect 248962 184170 249018 184226
rect 248838 184046 248894 184102
rect 248962 184046 249018 184102
rect 248838 183922 248894 183978
rect 248962 183922 249018 183978
rect 248838 166294 248894 166350
rect 248962 166294 249018 166350
rect 248838 166170 248894 166226
rect 248962 166170 249018 166226
rect 248838 166046 248894 166102
rect 248962 166046 249018 166102
rect 248838 165922 248894 165978
rect 248962 165922 249018 165978
rect 254994 298294 255050 298350
rect 255118 298294 255174 298350
rect 255242 298294 255298 298350
rect 255366 298294 255422 298350
rect 254994 298170 255050 298226
rect 255118 298170 255174 298226
rect 255242 298170 255298 298226
rect 255366 298170 255422 298226
rect 254994 298046 255050 298102
rect 255118 298046 255174 298102
rect 255242 298046 255298 298102
rect 255366 298046 255422 298102
rect 254994 297922 255050 297978
rect 255118 297922 255174 297978
rect 255242 297922 255298 297978
rect 255366 297922 255422 297978
rect 251274 274294 251330 274350
rect 251398 274294 251454 274350
rect 251522 274294 251578 274350
rect 251646 274294 251702 274350
rect 251274 274170 251330 274226
rect 251398 274170 251454 274226
rect 251522 274170 251578 274226
rect 251646 274170 251702 274226
rect 251274 274046 251330 274102
rect 251398 274046 251454 274102
rect 251522 274046 251578 274102
rect 251646 274046 251702 274102
rect 251274 273922 251330 273978
rect 251398 273922 251454 273978
rect 251522 273922 251578 273978
rect 251646 273922 251702 273978
rect 251274 256294 251330 256350
rect 251398 256294 251454 256350
rect 251522 256294 251578 256350
rect 251646 256294 251702 256350
rect 251274 256170 251330 256226
rect 251398 256170 251454 256226
rect 251522 256170 251578 256226
rect 251646 256170 251702 256226
rect 251274 256046 251330 256102
rect 251398 256046 251454 256102
rect 251522 256046 251578 256102
rect 251646 256046 251702 256102
rect 251274 255922 251330 255978
rect 251398 255922 251454 255978
rect 251522 255922 251578 255978
rect 251646 255922 251702 255978
rect 251274 238294 251330 238350
rect 251398 238294 251454 238350
rect 251522 238294 251578 238350
rect 251646 238294 251702 238350
rect 251274 238170 251330 238226
rect 251398 238170 251454 238226
rect 251522 238170 251578 238226
rect 251646 238170 251702 238226
rect 251274 238046 251330 238102
rect 251398 238046 251454 238102
rect 251522 238046 251578 238102
rect 251646 238046 251702 238102
rect 251274 237922 251330 237978
rect 251398 237922 251454 237978
rect 251522 237922 251578 237978
rect 251646 237922 251702 237978
rect 251274 220294 251330 220350
rect 251398 220294 251454 220350
rect 251522 220294 251578 220350
rect 251646 220294 251702 220350
rect 251274 220170 251330 220226
rect 251398 220170 251454 220226
rect 251522 220170 251578 220226
rect 251646 220170 251702 220226
rect 251274 220046 251330 220102
rect 251398 220046 251454 220102
rect 251522 220046 251578 220102
rect 251646 220046 251702 220102
rect 251274 219922 251330 219978
rect 251398 219922 251454 219978
rect 251522 219922 251578 219978
rect 251646 219922 251702 219978
rect 251274 202294 251330 202350
rect 251398 202294 251454 202350
rect 251522 202294 251578 202350
rect 251646 202294 251702 202350
rect 251274 202170 251330 202226
rect 251398 202170 251454 202226
rect 251522 202170 251578 202226
rect 251646 202170 251702 202226
rect 251274 202046 251330 202102
rect 251398 202046 251454 202102
rect 251522 202046 251578 202102
rect 251646 202046 251702 202102
rect 251274 201922 251330 201978
rect 251398 201922 251454 201978
rect 251522 201922 251578 201978
rect 251646 201922 251702 201978
rect 251274 184294 251330 184350
rect 251398 184294 251454 184350
rect 251522 184294 251578 184350
rect 251646 184294 251702 184350
rect 251274 184170 251330 184226
rect 251398 184170 251454 184226
rect 251522 184170 251578 184226
rect 251646 184170 251702 184226
rect 251274 184046 251330 184102
rect 251398 184046 251454 184102
rect 251522 184046 251578 184102
rect 251646 184046 251702 184102
rect 251274 183922 251330 183978
rect 251398 183922 251454 183978
rect 251522 183922 251578 183978
rect 251646 183922 251702 183978
rect 251274 166294 251330 166350
rect 251398 166294 251454 166350
rect 251522 166294 251578 166350
rect 251646 166294 251702 166350
rect 251274 166170 251330 166226
rect 251398 166170 251454 166226
rect 251522 166170 251578 166226
rect 251646 166170 251702 166226
rect 251274 166046 251330 166102
rect 251398 166046 251454 166102
rect 251522 166046 251578 166102
rect 251646 166046 251702 166102
rect 251274 165922 251330 165978
rect 251398 165922 251454 165978
rect 251522 165922 251578 165978
rect 251646 165922 251702 165978
rect 251274 148294 251330 148350
rect 251398 148294 251454 148350
rect 251522 148294 251578 148350
rect 251646 148294 251702 148350
rect 251274 148170 251330 148226
rect 251398 148170 251454 148226
rect 251522 148170 251578 148226
rect 251646 148170 251702 148226
rect 251274 148046 251330 148102
rect 251398 148046 251454 148102
rect 251522 148046 251578 148102
rect 251646 148046 251702 148102
rect 251274 147922 251330 147978
rect 251398 147922 251454 147978
rect 251522 147922 251578 147978
rect 251646 147922 251702 147978
rect 251274 130294 251330 130350
rect 251398 130294 251454 130350
rect 251522 130294 251578 130350
rect 251646 130294 251702 130350
rect 251274 130170 251330 130226
rect 251398 130170 251454 130226
rect 251522 130170 251578 130226
rect 251646 130170 251702 130226
rect 251274 130046 251330 130102
rect 251398 130046 251454 130102
rect 251522 130046 251578 130102
rect 251646 130046 251702 130102
rect 251274 129922 251330 129978
rect 251398 129922 251454 129978
rect 251522 129922 251578 129978
rect 251646 129922 251702 129978
rect 251274 112294 251330 112350
rect 251398 112294 251454 112350
rect 251522 112294 251578 112350
rect 251646 112294 251702 112350
rect 251274 112170 251330 112226
rect 251398 112170 251454 112226
rect 251522 112170 251578 112226
rect 251646 112170 251702 112226
rect 251274 112046 251330 112102
rect 251398 112046 251454 112102
rect 251522 112046 251578 112102
rect 251646 112046 251702 112102
rect 251274 111922 251330 111978
rect 251398 111922 251454 111978
rect 251522 111922 251578 111978
rect 251646 111922 251702 111978
rect 251274 94294 251330 94350
rect 251398 94294 251454 94350
rect 251522 94294 251578 94350
rect 251646 94294 251702 94350
rect 251274 94170 251330 94226
rect 251398 94170 251454 94226
rect 251522 94170 251578 94226
rect 251646 94170 251702 94226
rect 251274 94046 251330 94102
rect 251398 94046 251454 94102
rect 251522 94046 251578 94102
rect 251646 94046 251702 94102
rect 251274 93922 251330 93978
rect 251398 93922 251454 93978
rect 251522 93922 251578 93978
rect 251646 93922 251702 93978
rect 251274 76294 251330 76350
rect 251398 76294 251454 76350
rect 251522 76294 251578 76350
rect 251646 76294 251702 76350
rect 251274 76170 251330 76226
rect 251398 76170 251454 76226
rect 251522 76170 251578 76226
rect 251646 76170 251702 76226
rect 251274 76046 251330 76102
rect 251398 76046 251454 76102
rect 251522 76046 251578 76102
rect 251646 76046 251702 76102
rect 251274 75922 251330 75978
rect 251398 75922 251454 75978
rect 251522 75922 251578 75978
rect 251646 75922 251702 75978
rect 251274 58294 251330 58350
rect 251398 58294 251454 58350
rect 251522 58294 251578 58350
rect 251646 58294 251702 58350
rect 251274 58170 251330 58226
rect 251398 58170 251454 58226
rect 251522 58170 251578 58226
rect 251646 58170 251702 58226
rect 251274 58046 251330 58102
rect 251398 58046 251454 58102
rect 251522 58046 251578 58102
rect 251646 58046 251702 58102
rect 251274 57922 251330 57978
rect 251398 57922 251454 57978
rect 251522 57922 251578 57978
rect 251646 57922 251702 57978
rect 251274 40294 251330 40350
rect 251398 40294 251454 40350
rect 251522 40294 251578 40350
rect 251646 40294 251702 40350
rect 251274 40170 251330 40226
rect 251398 40170 251454 40226
rect 251522 40170 251578 40226
rect 251646 40170 251702 40226
rect 251274 40046 251330 40102
rect 251398 40046 251454 40102
rect 251522 40046 251578 40102
rect 251646 40046 251702 40102
rect 251274 39922 251330 39978
rect 251398 39922 251454 39978
rect 251522 39922 251578 39978
rect 251646 39922 251702 39978
rect 251274 22294 251330 22350
rect 251398 22294 251454 22350
rect 251522 22294 251578 22350
rect 251646 22294 251702 22350
rect 251274 22170 251330 22226
rect 251398 22170 251454 22226
rect 251522 22170 251578 22226
rect 251646 22170 251702 22226
rect 251274 22046 251330 22102
rect 251398 22046 251454 22102
rect 251522 22046 251578 22102
rect 251646 22046 251702 22102
rect 251274 21922 251330 21978
rect 251398 21922 251454 21978
rect 251522 21922 251578 21978
rect 251646 21922 251702 21978
rect 264198 298294 264254 298350
rect 264322 298294 264378 298350
rect 264198 298170 264254 298226
rect 264322 298170 264378 298226
rect 264198 298046 264254 298102
rect 264322 298046 264378 298102
rect 264198 297922 264254 297978
rect 264322 297922 264378 297978
rect 254994 280294 255050 280350
rect 255118 280294 255174 280350
rect 255242 280294 255298 280350
rect 255366 280294 255422 280350
rect 254994 280170 255050 280226
rect 255118 280170 255174 280226
rect 255242 280170 255298 280226
rect 255366 280170 255422 280226
rect 254994 280046 255050 280102
rect 255118 280046 255174 280102
rect 255242 280046 255298 280102
rect 255366 280046 255422 280102
rect 254994 279922 255050 279978
rect 255118 279922 255174 279978
rect 255242 279922 255298 279978
rect 255366 279922 255422 279978
rect 254994 262294 255050 262350
rect 255118 262294 255174 262350
rect 255242 262294 255298 262350
rect 255366 262294 255422 262350
rect 254994 262170 255050 262226
rect 255118 262170 255174 262226
rect 255242 262170 255298 262226
rect 255366 262170 255422 262226
rect 254994 262046 255050 262102
rect 255118 262046 255174 262102
rect 255242 262046 255298 262102
rect 255366 262046 255422 262102
rect 254994 261922 255050 261978
rect 255118 261922 255174 261978
rect 255242 261922 255298 261978
rect 255366 261922 255422 261978
rect 254994 244294 255050 244350
rect 255118 244294 255174 244350
rect 255242 244294 255298 244350
rect 255366 244294 255422 244350
rect 254994 244170 255050 244226
rect 255118 244170 255174 244226
rect 255242 244170 255298 244226
rect 255366 244170 255422 244226
rect 254994 244046 255050 244102
rect 255118 244046 255174 244102
rect 255242 244046 255298 244102
rect 255366 244046 255422 244102
rect 254994 243922 255050 243978
rect 255118 243922 255174 243978
rect 255242 243922 255298 243978
rect 255366 243922 255422 243978
rect 254994 226294 255050 226350
rect 255118 226294 255174 226350
rect 255242 226294 255298 226350
rect 255366 226294 255422 226350
rect 254994 226170 255050 226226
rect 255118 226170 255174 226226
rect 255242 226170 255298 226226
rect 255366 226170 255422 226226
rect 254994 226046 255050 226102
rect 255118 226046 255174 226102
rect 255242 226046 255298 226102
rect 255366 226046 255422 226102
rect 254994 225922 255050 225978
rect 255118 225922 255174 225978
rect 255242 225922 255298 225978
rect 255366 225922 255422 225978
rect 254994 208294 255050 208350
rect 255118 208294 255174 208350
rect 255242 208294 255298 208350
rect 255366 208294 255422 208350
rect 254994 208170 255050 208226
rect 255118 208170 255174 208226
rect 255242 208170 255298 208226
rect 255366 208170 255422 208226
rect 254994 208046 255050 208102
rect 255118 208046 255174 208102
rect 255242 208046 255298 208102
rect 255366 208046 255422 208102
rect 254994 207922 255050 207978
rect 255118 207922 255174 207978
rect 255242 207922 255298 207978
rect 255366 207922 255422 207978
rect 254994 190294 255050 190350
rect 255118 190294 255174 190350
rect 255242 190294 255298 190350
rect 255366 190294 255422 190350
rect 254994 190170 255050 190226
rect 255118 190170 255174 190226
rect 255242 190170 255298 190226
rect 255366 190170 255422 190226
rect 254994 190046 255050 190102
rect 255118 190046 255174 190102
rect 255242 190046 255298 190102
rect 255366 190046 255422 190102
rect 254994 189922 255050 189978
rect 255118 189922 255174 189978
rect 255242 189922 255298 189978
rect 255366 189922 255422 189978
rect 254994 172294 255050 172350
rect 255118 172294 255174 172350
rect 255242 172294 255298 172350
rect 255366 172294 255422 172350
rect 254994 172170 255050 172226
rect 255118 172170 255174 172226
rect 255242 172170 255298 172226
rect 255366 172170 255422 172226
rect 254994 172046 255050 172102
rect 255118 172046 255174 172102
rect 255242 172046 255298 172102
rect 255366 172046 255422 172102
rect 254994 171922 255050 171978
rect 255118 171922 255174 171978
rect 255242 171922 255298 171978
rect 255366 171922 255422 171978
rect 254994 154294 255050 154350
rect 255118 154294 255174 154350
rect 255242 154294 255298 154350
rect 255366 154294 255422 154350
rect 254994 154170 255050 154226
rect 255118 154170 255174 154226
rect 255242 154170 255298 154226
rect 255366 154170 255422 154226
rect 254994 154046 255050 154102
rect 255118 154046 255174 154102
rect 255242 154046 255298 154102
rect 255366 154046 255422 154102
rect 254994 153922 255050 153978
rect 255118 153922 255174 153978
rect 255242 153922 255298 153978
rect 255366 153922 255422 153978
rect 254994 136294 255050 136350
rect 255118 136294 255174 136350
rect 255242 136294 255298 136350
rect 255366 136294 255422 136350
rect 254994 136170 255050 136226
rect 255118 136170 255174 136226
rect 255242 136170 255298 136226
rect 255366 136170 255422 136226
rect 254994 136046 255050 136102
rect 255118 136046 255174 136102
rect 255242 136046 255298 136102
rect 255366 136046 255422 136102
rect 254994 135922 255050 135978
rect 255118 135922 255174 135978
rect 255242 135922 255298 135978
rect 255366 135922 255422 135978
rect 254994 118294 255050 118350
rect 255118 118294 255174 118350
rect 255242 118294 255298 118350
rect 255366 118294 255422 118350
rect 254994 118170 255050 118226
rect 255118 118170 255174 118226
rect 255242 118170 255298 118226
rect 255366 118170 255422 118226
rect 254994 118046 255050 118102
rect 255118 118046 255174 118102
rect 255242 118046 255298 118102
rect 255366 118046 255422 118102
rect 254994 117922 255050 117978
rect 255118 117922 255174 117978
rect 255242 117922 255298 117978
rect 255366 117922 255422 117978
rect 254994 100294 255050 100350
rect 255118 100294 255174 100350
rect 255242 100294 255298 100350
rect 255366 100294 255422 100350
rect 254994 100170 255050 100226
rect 255118 100170 255174 100226
rect 255242 100170 255298 100226
rect 255366 100170 255422 100226
rect 254994 100046 255050 100102
rect 255118 100046 255174 100102
rect 255242 100046 255298 100102
rect 255366 100046 255422 100102
rect 254994 99922 255050 99978
rect 255118 99922 255174 99978
rect 255242 99922 255298 99978
rect 255366 99922 255422 99978
rect 254994 82294 255050 82350
rect 255118 82294 255174 82350
rect 255242 82294 255298 82350
rect 255366 82294 255422 82350
rect 254994 82170 255050 82226
rect 255118 82170 255174 82226
rect 255242 82170 255298 82226
rect 255366 82170 255422 82226
rect 254994 82046 255050 82102
rect 255118 82046 255174 82102
rect 255242 82046 255298 82102
rect 255366 82046 255422 82102
rect 254994 81922 255050 81978
rect 255118 81922 255174 81978
rect 255242 81922 255298 81978
rect 255366 81922 255422 81978
rect 254994 64294 255050 64350
rect 255118 64294 255174 64350
rect 255242 64294 255298 64350
rect 255366 64294 255422 64350
rect 254994 64170 255050 64226
rect 255118 64170 255174 64226
rect 255242 64170 255298 64226
rect 255366 64170 255422 64226
rect 254994 64046 255050 64102
rect 255118 64046 255174 64102
rect 255242 64046 255298 64102
rect 255366 64046 255422 64102
rect 254994 63922 255050 63978
rect 255118 63922 255174 63978
rect 255242 63922 255298 63978
rect 255366 63922 255422 63978
rect 254994 46294 255050 46350
rect 255118 46294 255174 46350
rect 255242 46294 255298 46350
rect 255366 46294 255422 46350
rect 254994 46170 255050 46226
rect 255118 46170 255174 46226
rect 255242 46170 255298 46226
rect 255366 46170 255422 46226
rect 254994 46046 255050 46102
rect 255118 46046 255174 46102
rect 255242 46046 255298 46102
rect 255366 46046 255422 46102
rect 254994 45922 255050 45978
rect 255118 45922 255174 45978
rect 255242 45922 255298 45978
rect 255366 45922 255422 45978
rect 264198 190294 264254 190350
rect 264322 190294 264378 190350
rect 264198 190170 264254 190226
rect 264322 190170 264378 190226
rect 264198 190046 264254 190102
rect 264322 190046 264378 190102
rect 264198 189922 264254 189978
rect 264322 189922 264378 189978
rect 264198 172294 264254 172350
rect 264322 172294 264378 172350
rect 264198 172170 264254 172226
rect 264322 172170 264378 172226
rect 264198 172046 264254 172102
rect 264322 172046 264378 172102
rect 264198 171922 264254 171978
rect 264322 171922 264378 171978
rect 261130 130294 261186 130350
rect 261254 130294 261310 130350
rect 261378 130294 261434 130350
rect 261502 130294 261558 130350
rect 261130 130170 261186 130226
rect 261254 130170 261310 130226
rect 261378 130170 261434 130226
rect 261502 130170 261558 130226
rect 261130 130046 261186 130102
rect 261254 130046 261310 130102
rect 261378 130046 261434 130102
rect 261502 130046 261558 130102
rect 261130 129922 261186 129978
rect 261254 129922 261310 129978
rect 261378 129922 261434 129978
rect 261502 129922 261558 129978
rect 261930 118294 261986 118350
rect 262054 118294 262110 118350
rect 262178 118294 262234 118350
rect 262302 118294 262358 118350
rect 261930 118170 261986 118226
rect 262054 118170 262110 118226
rect 262178 118170 262234 118226
rect 262302 118170 262358 118226
rect 261930 118046 261986 118102
rect 262054 118046 262110 118102
rect 262178 118046 262234 118102
rect 262302 118046 262358 118102
rect 261930 117922 261986 117978
rect 262054 117922 262110 117978
rect 262178 117922 262234 117978
rect 262302 117922 262358 117978
rect 261130 112294 261186 112350
rect 261254 112294 261310 112350
rect 261378 112294 261434 112350
rect 261502 112294 261558 112350
rect 261130 112170 261186 112226
rect 261254 112170 261310 112226
rect 261378 112170 261434 112226
rect 261502 112170 261558 112226
rect 261130 112046 261186 112102
rect 261254 112046 261310 112102
rect 261378 112046 261434 112102
rect 261502 112046 261558 112102
rect 261130 111922 261186 111978
rect 261254 111922 261310 111978
rect 261378 111922 261434 111978
rect 261502 111922 261558 111978
rect 261930 100294 261986 100350
rect 262054 100294 262110 100350
rect 262178 100294 262234 100350
rect 262302 100294 262358 100350
rect 261930 100170 261986 100226
rect 262054 100170 262110 100226
rect 262178 100170 262234 100226
rect 262302 100170 262358 100226
rect 261930 100046 261986 100102
rect 262054 100046 262110 100102
rect 262178 100046 262234 100102
rect 262302 100046 262358 100102
rect 261930 99922 261986 99978
rect 262054 99922 262110 99978
rect 262178 99922 262234 99978
rect 262302 99922 262358 99978
rect 261130 94294 261186 94350
rect 261254 94294 261310 94350
rect 261378 94294 261434 94350
rect 261502 94294 261558 94350
rect 261130 94170 261186 94226
rect 261254 94170 261310 94226
rect 261378 94170 261434 94226
rect 261502 94170 261558 94226
rect 261130 94046 261186 94102
rect 261254 94046 261310 94102
rect 261378 94046 261434 94102
rect 261502 94046 261558 94102
rect 261130 93922 261186 93978
rect 261254 93922 261310 93978
rect 261378 93922 261434 93978
rect 261502 93922 261558 93978
rect 261930 82294 261986 82350
rect 262054 82294 262110 82350
rect 262178 82294 262234 82350
rect 262302 82294 262358 82350
rect 261930 82170 261986 82226
rect 262054 82170 262110 82226
rect 262178 82170 262234 82226
rect 262302 82170 262358 82226
rect 261930 82046 261986 82102
rect 262054 82046 262110 82102
rect 262178 82046 262234 82102
rect 262302 82046 262358 82102
rect 261930 81922 261986 81978
rect 262054 81922 262110 81978
rect 262178 81922 262234 81978
rect 262302 81922 262358 81978
rect 261130 76294 261186 76350
rect 261254 76294 261310 76350
rect 261378 76294 261434 76350
rect 261502 76294 261558 76350
rect 261130 76170 261186 76226
rect 261254 76170 261310 76226
rect 261378 76170 261434 76226
rect 261502 76170 261558 76226
rect 261130 76046 261186 76102
rect 261254 76046 261310 76102
rect 261378 76046 261434 76102
rect 261502 76046 261558 76102
rect 261130 75922 261186 75978
rect 261254 75922 261310 75978
rect 261378 75922 261434 75978
rect 261502 75922 261558 75978
rect 261930 64294 261986 64350
rect 262054 64294 262110 64350
rect 262178 64294 262234 64350
rect 262302 64294 262358 64350
rect 261930 64170 261986 64226
rect 262054 64170 262110 64226
rect 262178 64170 262234 64226
rect 262302 64170 262358 64226
rect 261930 64046 261986 64102
rect 262054 64046 262110 64102
rect 262178 64046 262234 64102
rect 262302 64046 262358 64102
rect 261930 63922 261986 63978
rect 262054 63922 262110 63978
rect 262178 63922 262234 63978
rect 262302 63922 262358 63978
rect 261130 58294 261186 58350
rect 261254 58294 261310 58350
rect 261378 58294 261434 58350
rect 261502 58294 261558 58350
rect 261130 58170 261186 58226
rect 261254 58170 261310 58226
rect 261378 58170 261434 58226
rect 261502 58170 261558 58226
rect 261130 58046 261186 58102
rect 261254 58046 261310 58102
rect 261378 58046 261434 58102
rect 261502 58046 261558 58102
rect 261130 57922 261186 57978
rect 261254 57922 261310 57978
rect 261378 57922 261434 57978
rect 261502 57922 261558 57978
rect 261930 46294 261986 46350
rect 262054 46294 262110 46350
rect 262178 46294 262234 46350
rect 262302 46294 262358 46350
rect 261930 46170 261986 46226
rect 262054 46170 262110 46226
rect 262178 46170 262234 46226
rect 262302 46170 262358 46226
rect 261930 46046 261986 46102
rect 262054 46046 262110 46102
rect 262178 46046 262234 46102
rect 262302 46046 262358 46102
rect 261930 45922 261986 45978
rect 262054 45922 262110 45978
rect 262178 45922 262234 45978
rect 262302 45922 262358 45978
rect 254994 28294 255050 28350
rect 255118 28294 255174 28350
rect 255242 28294 255298 28350
rect 255366 28294 255422 28350
rect 254994 28170 255050 28226
rect 255118 28170 255174 28226
rect 255242 28170 255298 28226
rect 255366 28170 255422 28226
rect 254994 28046 255050 28102
rect 255118 28046 255174 28102
rect 255242 28046 255298 28102
rect 255366 28046 255422 28102
rect 254994 27922 255050 27978
rect 255118 27922 255174 27978
rect 255242 27922 255298 27978
rect 255366 27922 255422 27978
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 276332 307502 276388 307558
rect 281372 427202 281428 427258
rect 281372 345662 281428 345718
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 285714 568294 285770 568350
rect 285838 568294 285894 568350
rect 285962 568294 286018 568350
rect 286086 568294 286142 568350
rect 285714 568170 285770 568226
rect 285838 568170 285894 568226
rect 285962 568170 286018 568226
rect 286086 568170 286142 568226
rect 285714 568046 285770 568102
rect 285838 568046 285894 568102
rect 285962 568046 286018 568102
rect 286086 568046 286142 568102
rect 285714 567922 285770 567978
rect 285838 567922 285894 567978
rect 285962 567922 286018 567978
rect 286086 567922 286142 567978
rect 285714 550294 285770 550350
rect 285838 550294 285894 550350
rect 285962 550294 286018 550350
rect 286086 550294 286142 550350
rect 285714 550170 285770 550226
rect 285838 550170 285894 550226
rect 285962 550170 286018 550226
rect 286086 550170 286142 550226
rect 285714 550046 285770 550102
rect 285838 550046 285894 550102
rect 285962 550046 286018 550102
rect 286086 550046 286142 550102
rect 285714 549922 285770 549978
rect 285838 549922 285894 549978
rect 285962 549922 286018 549978
rect 286086 549922 286142 549978
rect 285714 532294 285770 532350
rect 285838 532294 285894 532350
rect 285962 532294 286018 532350
rect 286086 532294 286142 532350
rect 285714 532170 285770 532226
rect 285838 532170 285894 532226
rect 285962 532170 286018 532226
rect 286086 532170 286142 532226
rect 285714 532046 285770 532102
rect 285838 532046 285894 532102
rect 285962 532046 286018 532102
rect 286086 532046 286142 532102
rect 285714 531922 285770 531978
rect 285838 531922 285894 531978
rect 285962 531922 286018 531978
rect 286086 531922 286142 531978
rect 285714 514294 285770 514350
rect 285838 514294 285894 514350
rect 285962 514294 286018 514350
rect 286086 514294 286142 514350
rect 285714 514170 285770 514226
rect 285838 514170 285894 514226
rect 285962 514170 286018 514226
rect 286086 514170 286142 514226
rect 285714 514046 285770 514102
rect 285838 514046 285894 514102
rect 285962 514046 286018 514102
rect 286086 514046 286142 514102
rect 285714 513922 285770 513978
rect 285838 513922 285894 513978
rect 285962 513922 286018 513978
rect 286086 513922 286142 513978
rect 285714 496294 285770 496350
rect 285838 496294 285894 496350
rect 285962 496294 286018 496350
rect 286086 496294 286142 496350
rect 285714 496170 285770 496226
rect 285838 496170 285894 496226
rect 285962 496170 286018 496226
rect 286086 496170 286142 496226
rect 285714 496046 285770 496102
rect 285838 496046 285894 496102
rect 285962 496046 286018 496102
rect 286086 496046 286142 496102
rect 285714 495922 285770 495978
rect 285838 495922 285894 495978
rect 285962 495922 286018 495978
rect 286086 495922 286142 495978
rect 285714 478294 285770 478350
rect 285838 478294 285894 478350
rect 285962 478294 286018 478350
rect 286086 478294 286142 478350
rect 285714 478170 285770 478226
rect 285838 478170 285894 478226
rect 285962 478170 286018 478226
rect 286086 478170 286142 478226
rect 285714 478046 285770 478102
rect 285838 478046 285894 478102
rect 285962 478046 286018 478102
rect 286086 478046 286142 478102
rect 285714 477922 285770 477978
rect 285838 477922 285894 477978
rect 285962 477922 286018 477978
rect 286086 477922 286142 477978
rect 285714 460294 285770 460350
rect 285838 460294 285894 460350
rect 285962 460294 286018 460350
rect 286086 460294 286142 460350
rect 285714 460170 285770 460226
rect 285838 460170 285894 460226
rect 285962 460170 286018 460226
rect 286086 460170 286142 460226
rect 285714 460046 285770 460102
rect 285838 460046 285894 460102
rect 285962 460046 286018 460102
rect 286086 460046 286142 460102
rect 285714 459922 285770 459978
rect 285838 459922 285894 459978
rect 285962 459922 286018 459978
rect 286086 459922 286142 459978
rect 285714 442294 285770 442350
rect 285838 442294 285894 442350
rect 285962 442294 286018 442350
rect 286086 442294 286142 442350
rect 285714 442170 285770 442226
rect 285838 442170 285894 442226
rect 285962 442170 286018 442226
rect 286086 442170 286142 442226
rect 285714 442046 285770 442102
rect 285838 442046 285894 442102
rect 285962 442046 286018 442102
rect 286086 442046 286142 442102
rect 285714 441922 285770 441978
rect 285838 441922 285894 441978
rect 285962 441922 286018 441978
rect 286086 441922 286142 441978
rect 284844 429362 284900 429418
rect 281994 418294 282050 418350
rect 282118 418294 282174 418350
rect 282242 418294 282298 418350
rect 282366 418294 282422 418350
rect 281994 418170 282050 418226
rect 282118 418170 282174 418226
rect 282242 418170 282298 418226
rect 282366 418170 282422 418226
rect 281994 418046 282050 418102
rect 282118 418046 282174 418102
rect 282242 418046 282298 418102
rect 282366 418046 282422 418102
rect 281994 417922 282050 417978
rect 282118 417922 282174 417978
rect 282242 417922 282298 417978
rect 282366 417922 282422 417978
rect 281994 400294 282050 400350
rect 282118 400294 282174 400350
rect 282242 400294 282298 400350
rect 282366 400294 282422 400350
rect 281994 400170 282050 400226
rect 282118 400170 282174 400226
rect 282242 400170 282298 400226
rect 282366 400170 282422 400226
rect 281994 400046 282050 400102
rect 282118 400046 282174 400102
rect 282242 400046 282298 400102
rect 282366 400046 282422 400102
rect 281994 399922 282050 399978
rect 282118 399922 282174 399978
rect 282242 399922 282298 399978
rect 282366 399922 282422 399978
rect 281994 382294 282050 382350
rect 282118 382294 282174 382350
rect 282242 382294 282298 382350
rect 282366 382294 282422 382350
rect 281994 382170 282050 382226
rect 282118 382170 282174 382226
rect 282242 382170 282298 382226
rect 282366 382170 282422 382226
rect 281994 382046 282050 382102
rect 282118 382046 282174 382102
rect 282242 382046 282298 382102
rect 282366 382046 282422 382102
rect 281994 381922 282050 381978
rect 282118 381922 282174 381978
rect 282242 381922 282298 381978
rect 282366 381922 282422 381978
rect 281994 364294 282050 364350
rect 282118 364294 282174 364350
rect 282242 364294 282298 364350
rect 282366 364294 282422 364350
rect 281994 364170 282050 364226
rect 282118 364170 282174 364226
rect 282242 364170 282298 364226
rect 282366 364170 282422 364226
rect 281994 364046 282050 364102
rect 282118 364046 282174 364102
rect 282242 364046 282298 364102
rect 282366 364046 282422 364102
rect 281994 363922 282050 363978
rect 282118 363922 282174 363978
rect 282242 363922 282298 363978
rect 282366 363922 282422 363978
rect 281994 346294 282050 346350
rect 282118 346294 282174 346350
rect 282242 346294 282298 346350
rect 282366 346294 282422 346350
rect 281994 346170 282050 346226
rect 282118 346170 282174 346226
rect 282242 346170 282298 346226
rect 282366 346170 282422 346226
rect 281994 346046 282050 346102
rect 282118 346046 282174 346102
rect 282242 346046 282298 346102
rect 282366 346046 282422 346102
rect 281994 345922 282050 345978
rect 282118 345922 282174 345978
rect 282242 345922 282298 345978
rect 282366 345922 282422 345978
rect 279692 337562 279748 337618
rect 283052 423422 283108 423478
rect 283052 330902 283108 330958
rect 281994 328294 282050 328350
rect 282118 328294 282174 328350
rect 282242 328294 282298 328350
rect 282366 328294 282422 328350
rect 281994 328170 282050 328226
rect 282118 328170 282174 328226
rect 282242 328170 282298 328226
rect 282366 328170 282422 328226
rect 281994 328046 282050 328102
rect 282118 328046 282174 328102
rect 282242 328046 282298 328102
rect 282366 328046 282422 328102
rect 281994 327922 282050 327978
rect 282118 327922 282174 327978
rect 282242 327922 282298 327978
rect 282366 327922 282422 327978
rect 281372 312542 281428 312598
rect 281994 310294 282050 310350
rect 282118 310294 282174 310350
rect 282242 310294 282298 310350
rect 282366 310294 282422 310350
rect 281994 310170 282050 310226
rect 282118 310170 282174 310226
rect 282242 310170 282298 310226
rect 282366 310170 282422 310226
rect 281994 310046 282050 310102
rect 282118 310046 282174 310102
rect 282242 310046 282298 310102
rect 282366 310046 282422 310102
rect 281994 309922 282050 309978
rect 282118 309922 282174 309978
rect 282242 309922 282298 309978
rect 282366 309922 282422 309978
rect 281994 292294 282050 292350
rect 282118 292294 282174 292350
rect 282242 292294 282298 292350
rect 282366 292294 282422 292350
rect 281994 292170 282050 292226
rect 282118 292170 282174 292226
rect 282242 292170 282298 292226
rect 282366 292170 282422 292226
rect 281994 292046 282050 292102
rect 282118 292046 282174 292102
rect 282242 292046 282298 292102
rect 282366 292046 282422 292102
rect 283052 321002 283108 321058
rect 281994 291922 282050 291978
rect 282118 291922 282174 291978
rect 282242 291922 282298 291978
rect 282366 291922 282422 291978
rect 281994 274294 282050 274350
rect 282118 274294 282174 274350
rect 282242 274294 282298 274350
rect 282366 274294 282422 274350
rect 281994 274170 282050 274226
rect 282118 274170 282174 274226
rect 282242 274170 282298 274226
rect 282366 274170 282422 274226
rect 281994 274046 282050 274102
rect 282118 274046 282174 274102
rect 282242 274046 282298 274102
rect 282366 274046 282422 274102
rect 281994 273922 282050 273978
rect 282118 273922 282174 273978
rect 282242 273922 282298 273978
rect 282366 273922 282422 273978
rect 281994 256294 282050 256350
rect 282118 256294 282174 256350
rect 282242 256294 282298 256350
rect 282366 256294 282422 256350
rect 281994 256170 282050 256226
rect 282118 256170 282174 256226
rect 282242 256170 282298 256226
rect 282366 256170 282422 256226
rect 281994 256046 282050 256102
rect 282118 256046 282174 256102
rect 282242 256046 282298 256102
rect 282366 256046 282422 256102
rect 281994 255922 282050 255978
rect 282118 255922 282174 255978
rect 282242 255922 282298 255978
rect 282366 255922 282422 255978
rect 281994 238294 282050 238350
rect 282118 238294 282174 238350
rect 282242 238294 282298 238350
rect 282366 238294 282422 238350
rect 281994 238170 282050 238226
rect 282118 238170 282174 238226
rect 282242 238170 282298 238226
rect 282366 238170 282422 238226
rect 281994 238046 282050 238102
rect 282118 238046 282174 238102
rect 282242 238046 282298 238102
rect 282366 238046 282422 238102
rect 281994 237922 282050 237978
rect 282118 237922 282174 237978
rect 282242 237922 282298 237978
rect 282366 237922 282422 237978
rect 281994 220294 282050 220350
rect 282118 220294 282174 220350
rect 282242 220294 282298 220350
rect 282366 220294 282422 220350
rect 281994 220170 282050 220226
rect 282118 220170 282174 220226
rect 282242 220170 282298 220226
rect 282366 220170 282422 220226
rect 281994 220046 282050 220102
rect 282118 220046 282174 220102
rect 282242 220046 282298 220102
rect 282366 220046 282422 220102
rect 281994 219922 282050 219978
rect 282118 219922 282174 219978
rect 282242 219922 282298 219978
rect 282366 219922 282422 219978
rect 281994 202294 282050 202350
rect 282118 202294 282174 202350
rect 282242 202294 282298 202350
rect 282366 202294 282422 202350
rect 281994 202170 282050 202226
rect 282118 202170 282174 202226
rect 282242 202170 282298 202226
rect 282366 202170 282422 202226
rect 281994 202046 282050 202102
rect 282118 202046 282174 202102
rect 282242 202046 282298 202102
rect 282366 202046 282422 202102
rect 281994 201922 282050 201978
rect 282118 201922 282174 201978
rect 282242 201922 282298 201978
rect 282366 201922 282422 201978
rect 281994 184294 282050 184350
rect 282118 184294 282174 184350
rect 282242 184294 282298 184350
rect 282366 184294 282422 184350
rect 281994 184170 282050 184226
rect 282118 184170 282174 184226
rect 282242 184170 282298 184226
rect 282366 184170 282422 184226
rect 281994 184046 282050 184102
rect 282118 184046 282174 184102
rect 282242 184046 282298 184102
rect 282366 184046 282422 184102
rect 281994 183922 282050 183978
rect 282118 183922 282174 183978
rect 282242 183922 282298 183978
rect 282366 183922 282422 183978
rect 281994 166294 282050 166350
rect 282118 166294 282174 166350
rect 282242 166294 282298 166350
rect 282366 166294 282422 166350
rect 281994 166170 282050 166226
rect 282118 166170 282174 166226
rect 282242 166170 282298 166226
rect 282366 166170 282422 166226
rect 281994 166046 282050 166102
rect 282118 166046 282174 166102
rect 282242 166046 282298 166102
rect 282366 166046 282422 166102
rect 281994 165922 282050 165978
rect 282118 165922 282174 165978
rect 282242 165922 282298 165978
rect 282366 165922 282422 165978
rect 281994 148294 282050 148350
rect 282118 148294 282174 148350
rect 282242 148294 282298 148350
rect 282366 148294 282422 148350
rect 281994 148170 282050 148226
rect 282118 148170 282174 148226
rect 282242 148170 282298 148226
rect 282366 148170 282422 148226
rect 281994 148046 282050 148102
rect 282118 148046 282174 148102
rect 282242 148046 282298 148102
rect 282366 148046 282422 148102
rect 281994 147922 282050 147978
rect 282118 147922 282174 147978
rect 282242 147922 282298 147978
rect 282366 147922 282422 147978
rect 281994 130294 282050 130350
rect 282118 130294 282174 130350
rect 282242 130294 282298 130350
rect 282366 130294 282422 130350
rect 281994 130170 282050 130226
rect 282118 130170 282174 130226
rect 282242 130170 282298 130226
rect 282366 130170 282422 130226
rect 281994 130046 282050 130102
rect 282118 130046 282174 130102
rect 282242 130046 282298 130102
rect 282366 130046 282422 130102
rect 281994 129922 282050 129978
rect 282118 129922 282174 129978
rect 282242 129922 282298 129978
rect 282366 129922 282422 129978
rect 281994 112294 282050 112350
rect 282118 112294 282174 112350
rect 282242 112294 282298 112350
rect 282366 112294 282422 112350
rect 281994 112170 282050 112226
rect 282118 112170 282174 112226
rect 282242 112170 282298 112226
rect 282366 112170 282422 112226
rect 281994 112046 282050 112102
rect 282118 112046 282174 112102
rect 282242 112046 282298 112102
rect 282366 112046 282422 112102
rect 281994 111922 282050 111978
rect 282118 111922 282174 111978
rect 282242 111922 282298 111978
rect 282366 111922 282422 111978
rect 281994 94294 282050 94350
rect 282118 94294 282174 94350
rect 282242 94294 282298 94350
rect 282366 94294 282422 94350
rect 281994 94170 282050 94226
rect 282118 94170 282174 94226
rect 282242 94170 282298 94226
rect 282366 94170 282422 94226
rect 281994 94046 282050 94102
rect 282118 94046 282174 94102
rect 282242 94046 282298 94102
rect 282366 94046 282422 94102
rect 281994 93922 282050 93978
rect 282118 93922 282174 93978
rect 282242 93922 282298 93978
rect 282366 93922 282422 93978
rect 281994 76294 282050 76350
rect 282118 76294 282174 76350
rect 282242 76294 282298 76350
rect 282366 76294 282422 76350
rect 281994 76170 282050 76226
rect 282118 76170 282174 76226
rect 282242 76170 282298 76226
rect 282366 76170 282422 76226
rect 281994 76046 282050 76102
rect 282118 76046 282174 76102
rect 282242 76046 282298 76102
rect 282366 76046 282422 76102
rect 281994 75922 282050 75978
rect 282118 75922 282174 75978
rect 282242 75922 282298 75978
rect 282366 75922 282422 75978
rect 281994 58294 282050 58350
rect 282118 58294 282174 58350
rect 282242 58294 282298 58350
rect 282366 58294 282422 58350
rect 281994 58170 282050 58226
rect 282118 58170 282174 58226
rect 282242 58170 282298 58226
rect 282366 58170 282422 58226
rect 281994 58046 282050 58102
rect 282118 58046 282174 58102
rect 282242 58046 282298 58102
rect 282366 58046 282422 58102
rect 281994 57922 282050 57978
rect 282118 57922 282174 57978
rect 282242 57922 282298 57978
rect 282366 57922 282422 57978
rect 281994 40294 282050 40350
rect 282118 40294 282174 40350
rect 282242 40294 282298 40350
rect 282366 40294 282422 40350
rect 281994 40170 282050 40226
rect 282118 40170 282174 40226
rect 282242 40170 282298 40226
rect 282366 40170 282422 40226
rect 281994 40046 282050 40102
rect 282118 40046 282174 40102
rect 282242 40046 282298 40102
rect 282366 40046 282422 40102
rect 281994 39922 282050 39978
rect 282118 39922 282174 39978
rect 282242 39922 282298 39978
rect 282366 39922 282422 39978
rect 281994 22294 282050 22350
rect 282118 22294 282174 22350
rect 282242 22294 282298 22350
rect 282366 22294 282422 22350
rect 281994 22170 282050 22226
rect 282118 22170 282174 22226
rect 282242 22170 282298 22226
rect 282366 22170 282422 22226
rect 281994 22046 282050 22102
rect 282118 22046 282174 22102
rect 282242 22046 282298 22102
rect 282366 22046 282422 22102
rect 281994 21922 282050 21978
rect 282118 21922 282174 21978
rect 282242 21922 282298 21978
rect 282366 21922 282422 21978
rect 284956 345302 285012 345358
rect 288092 589742 288148 589798
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 312714 562294 312770 562350
rect 312838 562294 312894 562350
rect 312962 562294 313018 562350
rect 313086 562294 313142 562350
rect 312714 562170 312770 562226
rect 312838 562170 312894 562226
rect 312962 562170 313018 562226
rect 313086 562170 313142 562226
rect 312714 562046 312770 562102
rect 312838 562046 312894 562102
rect 312962 562046 313018 562102
rect 313086 562046 313142 562102
rect 312714 561922 312770 561978
rect 312838 561922 312894 561978
rect 312962 561922 313018 561978
rect 313086 561922 313142 561978
rect 300524 521724 300580 521758
rect 300524 521702 300580 521724
rect 300636 520268 300692 520318
rect 300636 520262 300692 520268
rect 300524 516852 300580 516898
rect 300524 516842 300580 516852
rect 300636 513604 300692 513658
rect 300636 513602 300692 513604
rect 301868 521702 301924 521758
rect 301756 520262 301812 520318
rect 301644 516842 301700 516898
rect 301532 513602 301588 513658
rect 303324 488042 303380 488098
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 316434 568294 316490 568350
rect 316558 568294 316614 568350
rect 316682 568294 316738 568350
rect 316806 568294 316862 568350
rect 316434 568170 316490 568226
rect 316558 568170 316614 568226
rect 316682 568170 316738 568226
rect 316806 568170 316862 568226
rect 316434 568046 316490 568102
rect 316558 568046 316614 568102
rect 316682 568046 316738 568102
rect 316806 568046 316862 568102
rect 316434 567922 316490 567978
rect 316558 567922 316614 567978
rect 316682 567922 316738 567978
rect 316806 567922 316862 567978
rect 316434 550294 316490 550350
rect 316558 550294 316614 550350
rect 316682 550294 316738 550350
rect 316806 550294 316862 550350
rect 316434 550170 316490 550226
rect 316558 550170 316614 550226
rect 316682 550170 316738 550226
rect 316806 550170 316862 550226
rect 316434 550046 316490 550102
rect 316558 550046 316614 550102
rect 316682 550046 316738 550102
rect 316806 550046 316862 550102
rect 316434 549922 316490 549978
rect 316558 549922 316614 549978
rect 316682 549922 316738 549978
rect 316806 549922 316862 549978
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 343434 562294 343490 562350
rect 343558 562294 343614 562350
rect 343682 562294 343738 562350
rect 343806 562294 343862 562350
rect 343434 562170 343490 562226
rect 343558 562170 343614 562226
rect 343682 562170 343738 562226
rect 343806 562170 343862 562226
rect 343434 562046 343490 562102
rect 343558 562046 343614 562102
rect 343682 562046 343738 562102
rect 343806 562046 343862 562102
rect 343434 561922 343490 561978
rect 343558 561922 343614 561978
rect 343682 561922 343738 561978
rect 343806 561922 343862 561978
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 347154 568294 347210 568350
rect 347278 568294 347334 568350
rect 347402 568294 347458 568350
rect 347526 568294 347582 568350
rect 347154 568170 347210 568226
rect 347278 568170 347334 568226
rect 347402 568170 347458 568226
rect 347526 568170 347582 568226
rect 347154 568046 347210 568102
rect 347278 568046 347334 568102
rect 347402 568046 347458 568102
rect 347526 568046 347582 568102
rect 347154 567922 347210 567978
rect 347278 567922 347334 567978
rect 347402 567922 347458 567978
rect 347526 567922 347582 567978
rect 347154 550294 347210 550350
rect 347278 550294 347334 550350
rect 347402 550294 347458 550350
rect 347526 550294 347582 550350
rect 347154 550170 347210 550226
rect 347278 550170 347334 550226
rect 347402 550170 347458 550226
rect 347526 550170 347582 550226
rect 347154 550046 347210 550102
rect 347278 550046 347334 550102
rect 347402 550046 347458 550102
rect 347526 550046 347582 550102
rect 347154 549922 347210 549978
rect 347278 549922 347334 549978
rect 347402 549922 347458 549978
rect 347526 549922 347582 549978
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 374154 562294 374210 562350
rect 374278 562294 374334 562350
rect 374402 562294 374458 562350
rect 374526 562294 374582 562350
rect 374154 562170 374210 562226
rect 374278 562170 374334 562226
rect 374402 562170 374458 562226
rect 374526 562170 374582 562226
rect 374154 562046 374210 562102
rect 374278 562046 374334 562102
rect 374402 562046 374458 562102
rect 374526 562046 374582 562102
rect 374154 561922 374210 561978
rect 374278 561922 374334 561978
rect 374402 561922 374458 561978
rect 374526 561922 374582 561978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 377874 568294 377930 568350
rect 377998 568294 378054 568350
rect 378122 568294 378178 568350
rect 378246 568294 378302 568350
rect 377874 568170 377930 568226
rect 377998 568170 378054 568226
rect 378122 568170 378178 568226
rect 378246 568170 378302 568226
rect 377874 568046 377930 568102
rect 377998 568046 378054 568102
rect 378122 568046 378178 568102
rect 378246 568046 378302 568102
rect 377874 567922 377930 567978
rect 377998 567922 378054 567978
rect 378122 567922 378178 567978
rect 378246 567922 378302 567978
rect 377874 550294 377930 550350
rect 377998 550294 378054 550350
rect 378122 550294 378178 550350
rect 378246 550294 378302 550350
rect 377874 550170 377930 550226
rect 377998 550170 378054 550226
rect 378122 550170 378178 550226
rect 378246 550170 378302 550226
rect 377874 550046 377930 550102
rect 377998 550046 378054 550102
rect 378122 550046 378178 550102
rect 378246 550046 378302 550102
rect 377874 549922 377930 549978
rect 377998 549922 378054 549978
rect 378122 549922 378178 549978
rect 378246 549922 378302 549978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 404874 562294 404930 562350
rect 404998 562294 405054 562350
rect 405122 562294 405178 562350
rect 405246 562294 405302 562350
rect 404874 562170 404930 562226
rect 404998 562170 405054 562226
rect 405122 562170 405178 562226
rect 405246 562170 405302 562226
rect 404874 562046 404930 562102
rect 404998 562046 405054 562102
rect 405122 562046 405178 562102
rect 405246 562046 405302 562102
rect 404874 561922 404930 561978
rect 404998 561922 405054 561978
rect 405122 561922 405178 561978
rect 405246 561922 405302 561978
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 408594 568294 408650 568350
rect 408718 568294 408774 568350
rect 408842 568294 408898 568350
rect 408966 568294 409022 568350
rect 408594 568170 408650 568226
rect 408718 568170 408774 568226
rect 408842 568170 408898 568226
rect 408966 568170 409022 568226
rect 408594 568046 408650 568102
rect 408718 568046 408774 568102
rect 408842 568046 408898 568102
rect 408966 568046 409022 568102
rect 408594 567922 408650 567978
rect 408718 567922 408774 567978
rect 408842 567922 408898 567978
rect 408966 567922 409022 567978
rect 408594 550294 408650 550350
rect 408718 550294 408774 550350
rect 408842 550294 408898 550350
rect 408966 550294 409022 550350
rect 408594 550170 408650 550226
rect 408718 550170 408774 550226
rect 408842 550170 408898 550226
rect 408966 550170 409022 550226
rect 408594 550046 408650 550102
rect 408718 550046 408774 550102
rect 408842 550046 408898 550102
rect 408966 550046 409022 550102
rect 408594 549922 408650 549978
rect 408718 549922 408774 549978
rect 408842 549922 408898 549978
rect 408966 549922 409022 549978
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 435594 562294 435650 562350
rect 435718 562294 435774 562350
rect 435842 562294 435898 562350
rect 435966 562294 436022 562350
rect 435594 562170 435650 562226
rect 435718 562170 435774 562226
rect 435842 562170 435898 562226
rect 435966 562170 436022 562226
rect 435594 562046 435650 562102
rect 435718 562046 435774 562102
rect 435842 562046 435898 562102
rect 435966 562046 436022 562102
rect 435594 561922 435650 561978
rect 435718 561922 435774 561978
rect 435842 561922 435898 561978
rect 435966 561922 436022 561978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 439314 568294 439370 568350
rect 439438 568294 439494 568350
rect 439562 568294 439618 568350
rect 439686 568294 439742 568350
rect 439314 568170 439370 568226
rect 439438 568170 439494 568226
rect 439562 568170 439618 568226
rect 439686 568170 439742 568226
rect 439314 568046 439370 568102
rect 439438 568046 439494 568102
rect 439562 568046 439618 568102
rect 439686 568046 439742 568102
rect 439314 567922 439370 567978
rect 439438 567922 439494 567978
rect 439562 567922 439618 567978
rect 439686 567922 439742 567978
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 466314 562294 466370 562350
rect 466438 562294 466494 562350
rect 466562 562294 466618 562350
rect 466686 562294 466742 562350
rect 466314 562170 466370 562226
rect 466438 562170 466494 562226
rect 466562 562170 466618 562226
rect 466686 562170 466742 562226
rect 466314 562046 466370 562102
rect 466438 562046 466494 562102
rect 466562 562046 466618 562102
rect 466686 562046 466742 562102
rect 466314 561922 466370 561978
rect 466438 561922 466494 561978
rect 466562 561922 466618 561978
rect 466686 561922 466742 561978
rect 459452 557882 459508 557938
rect 439314 550294 439370 550350
rect 439438 550294 439494 550350
rect 439562 550294 439618 550350
rect 439686 550294 439742 550350
rect 439314 550170 439370 550226
rect 439438 550170 439494 550226
rect 439562 550170 439618 550226
rect 439686 550170 439742 550226
rect 439314 550046 439370 550102
rect 439438 550046 439494 550102
rect 439562 550046 439618 550102
rect 439686 550046 439742 550102
rect 439314 549922 439370 549978
rect 439438 549922 439494 549978
rect 439562 549922 439618 549978
rect 439686 549922 439742 549978
rect 452732 551222 452788 551278
rect 304518 544294 304574 544350
rect 304642 544294 304698 544350
rect 304518 544170 304574 544226
rect 304642 544170 304698 544226
rect 304518 544046 304574 544102
rect 304642 544046 304698 544102
rect 304518 543922 304574 543978
rect 304642 543922 304698 543978
rect 335238 544294 335294 544350
rect 335362 544294 335418 544350
rect 335238 544170 335294 544226
rect 335362 544170 335418 544226
rect 335238 544046 335294 544102
rect 335362 544046 335418 544102
rect 335238 543922 335294 543978
rect 335362 543922 335418 543978
rect 365958 544294 366014 544350
rect 366082 544294 366138 544350
rect 365958 544170 366014 544226
rect 366082 544170 366138 544226
rect 365958 544046 366014 544102
rect 366082 544046 366138 544102
rect 365958 543922 366014 543978
rect 366082 543922 366138 543978
rect 396678 544294 396734 544350
rect 396802 544294 396858 544350
rect 396678 544170 396734 544226
rect 396802 544170 396858 544226
rect 396678 544046 396734 544102
rect 396802 544046 396858 544102
rect 396678 543922 396734 543978
rect 396802 543922 396858 543978
rect 427398 544294 427454 544350
rect 427522 544294 427578 544350
rect 427398 544170 427454 544226
rect 427522 544170 427578 544226
rect 427398 544046 427454 544102
rect 427522 544046 427578 544102
rect 427398 543922 427454 543978
rect 427522 543922 427578 543978
rect 319878 532294 319934 532350
rect 320002 532294 320058 532350
rect 319878 532170 319934 532226
rect 320002 532170 320058 532226
rect 319878 532046 319934 532102
rect 320002 532046 320058 532102
rect 319878 531922 319934 531978
rect 320002 531922 320058 531978
rect 350598 532294 350654 532350
rect 350722 532294 350778 532350
rect 350598 532170 350654 532226
rect 350722 532170 350778 532226
rect 350598 532046 350654 532102
rect 350722 532046 350778 532102
rect 350598 531922 350654 531978
rect 350722 531922 350778 531978
rect 381318 532294 381374 532350
rect 381442 532294 381498 532350
rect 381318 532170 381374 532226
rect 381442 532170 381498 532226
rect 381318 532046 381374 532102
rect 381442 532046 381498 532102
rect 381318 531922 381374 531978
rect 381442 531922 381498 531978
rect 412038 532294 412094 532350
rect 412162 532294 412218 532350
rect 412038 532170 412094 532226
rect 412162 532170 412218 532226
rect 412038 532046 412094 532102
rect 412162 532046 412218 532102
rect 412038 531922 412094 531978
rect 412162 531922 412218 531978
rect 442758 532294 442814 532350
rect 442882 532294 442938 532350
rect 442758 532170 442814 532226
rect 442882 532170 442938 532226
rect 442758 532046 442814 532102
rect 442882 532046 442938 532102
rect 442758 531922 442814 531978
rect 442882 531922 442938 531978
rect 304518 526294 304574 526350
rect 304642 526294 304698 526350
rect 304518 526170 304574 526226
rect 304642 526170 304698 526226
rect 304518 526046 304574 526102
rect 304642 526046 304698 526102
rect 304518 525922 304574 525978
rect 304642 525922 304698 525978
rect 335238 526294 335294 526350
rect 335362 526294 335418 526350
rect 335238 526170 335294 526226
rect 335362 526170 335418 526226
rect 335238 526046 335294 526102
rect 335362 526046 335418 526102
rect 335238 525922 335294 525978
rect 335362 525922 335418 525978
rect 365958 526294 366014 526350
rect 366082 526294 366138 526350
rect 365958 526170 366014 526226
rect 366082 526170 366138 526226
rect 365958 526046 366014 526102
rect 366082 526046 366138 526102
rect 365958 525922 366014 525978
rect 366082 525922 366138 525978
rect 396678 526294 396734 526350
rect 396802 526294 396858 526350
rect 396678 526170 396734 526226
rect 396802 526170 396858 526226
rect 396678 526046 396734 526102
rect 396802 526046 396858 526102
rect 396678 525922 396734 525978
rect 396802 525922 396858 525978
rect 427398 526294 427454 526350
rect 427522 526294 427578 526350
rect 427398 526170 427454 526226
rect 427522 526170 427578 526226
rect 427398 526046 427454 526102
rect 427522 526046 427578 526102
rect 427398 525922 427454 525978
rect 427522 525922 427578 525978
rect 319878 514294 319934 514350
rect 320002 514294 320058 514350
rect 319878 514170 319934 514226
rect 320002 514170 320058 514226
rect 319878 514046 319934 514102
rect 320002 514046 320058 514102
rect 319878 513922 319934 513978
rect 320002 513922 320058 513978
rect 350598 514294 350654 514350
rect 350722 514294 350778 514350
rect 350598 514170 350654 514226
rect 350722 514170 350778 514226
rect 350598 514046 350654 514102
rect 350722 514046 350778 514102
rect 350598 513922 350654 513978
rect 350722 513922 350778 513978
rect 381318 514294 381374 514350
rect 381442 514294 381498 514350
rect 381318 514170 381374 514226
rect 381442 514170 381498 514226
rect 381318 514046 381374 514102
rect 381442 514046 381498 514102
rect 381318 513922 381374 513978
rect 381442 513922 381498 513978
rect 412038 514294 412094 514350
rect 412162 514294 412218 514350
rect 412038 514170 412094 514226
rect 412162 514170 412218 514226
rect 412038 514046 412094 514102
rect 412162 514046 412218 514102
rect 412038 513922 412094 513978
rect 412162 513922 412218 513978
rect 442758 514294 442814 514350
rect 442882 514294 442938 514350
rect 442758 514170 442814 514226
rect 442882 514170 442938 514226
rect 442758 514046 442814 514102
rect 442882 514046 442938 514102
rect 442758 513922 442814 513978
rect 442882 513922 442938 513978
rect 304518 508294 304574 508350
rect 304642 508294 304698 508350
rect 304518 508170 304574 508226
rect 304642 508170 304698 508226
rect 304518 508046 304574 508102
rect 304642 508046 304698 508102
rect 304518 507922 304574 507978
rect 304642 507922 304698 507978
rect 335238 508294 335294 508350
rect 335362 508294 335418 508350
rect 335238 508170 335294 508226
rect 335362 508170 335418 508226
rect 335238 508046 335294 508102
rect 335362 508046 335418 508102
rect 335238 507922 335294 507978
rect 335362 507922 335418 507978
rect 365958 508294 366014 508350
rect 366082 508294 366138 508350
rect 365958 508170 366014 508226
rect 366082 508170 366138 508226
rect 365958 508046 366014 508102
rect 366082 508046 366138 508102
rect 365958 507922 366014 507978
rect 366082 507922 366138 507978
rect 396678 508294 396734 508350
rect 396802 508294 396858 508350
rect 396678 508170 396734 508226
rect 396802 508170 396858 508226
rect 396678 508046 396734 508102
rect 396802 508046 396858 508102
rect 396678 507922 396734 507978
rect 396802 507922 396858 507978
rect 427398 508294 427454 508350
rect 427522 508294 427578 508350
rect 427398 508170 427454 508226
rect 427522 508170 427578 508226
rect 427398 508046 427454 508102
rect 427522 508046 427578 508102
rect 427398 507922 427454 507978
rect 427522 507922 427578 507978
rect 446012 499742 446068 499798
rect 319878 496294 319934 496350
rect 320002 496294 320058 496350
rect 319878 496170 319934 496226
rect 320002 496170 320058 496226
rect 319878 496046 319934 496102
rect 320002 496046 320058 496102
rect 319878 495922 319934 495978
rect 320002 495922 320058 495978
rect 350598 496294 350654 496350
rect 350722 496294 350778 496350
rect 350598 496170 350654 496226
rect 350722 496170 350778 496226
rect 350598 496046 350654 496102
rect 350722 496046 350778 496102
rect 350598 495922 350654 495978
rect 350722 495922 350778 495978
rect 381318 496294 381374 496350
rect 381442 496294 381498 496350
rect 381318 496170 381374 496226
rect 381442 496170 381498 496226
rect 381318 496046 381374 496102
rect 381442 496046 381498 496102
rect 381318 495922 381374 495978
rect 381442 495922 381498 495978
rect 412038 496294 412094 496350
rect 412162 496294 412218 496350
rect 412038 496170 412094 496226
rect 412162 496170 412218 496226
rect 412038 496046 412094 496102
rect 412162 496046 412218 496102
rect 412038 495922 412094 495978
rect 412162 495922 412218 495978
rect 442758 496294 442814 496350
rect 442882 496294 442938 496350
rect 442758 496170 442814 496226
rect 442882 496170 442938 496226
rect 442758 496046 442814 496102
rect 442882 496046 442938 496102
rect 442758 495922 442814 495978
rect 442882 495922 442938 495978
rect 304518 490294 304574 490350
rect 304642 490294 304698 490350
rect 304518 490170 304574 490226
rect 304642 490170 304698 490226
rect 304518 490046 304574 490102
rect 304642 490046 304698 490102
rect 304518 489922 304574 489978
rect 304642 489922 304698 489978
rect 335238 490294 335294 490350
rect 335362 490294 335418 490350
rect 335238 490170 335294 490226
rect 335362 490170 335418 490226
rect 335238 490046 335294 490102
rect 335362 490046 335418 490102
rect 335238 489922 335294 489978
rect 335362 489922 335418 489978
rect 365958 490294 366014 490350
rect 366082 490294 366138 490350
rect 365958 490170 366014 490226
rect 366082 490170 366138 490226
rect 365958 490046 366014 490102
rect 366082 490046 366138 490102
rect 365958 489922 366014 489978
rect 366082 489922 366138 489978
rect 396678 490294 396734 490350
rect 396802 490294 396858 490350
rect 396678 490170 396734 490226
rect 396802 490170 396858 490226
rect 396678 490046 396734 490102
rect 396802 490046 396858 490102
rect 396678 489922 396734 489978
rect 396802 489922 396858 489978
rect 427398 490294 427454 490350
rect 427522 490294 427578 490350
rect 427398 490170 427454 490226
rect 427522 490170 427578 490226
rect 427398 490046 427454 490102
rect 427522 490046 427578 490102
rect 427398 489922 427454 489978
rect 427522 489922 427578 489978
rect 303436 479582 303492 479638
rect 319878 478294 319934 478350
rect 320002 478294 320058 478350
rect 319878 478170 319934 478226
rect 320002 478170 320058 478226
rect 319878 478046 319934 478102
rect 320002 478046 320058 478102
rect 319878 477922 319934 477978
rect 320002 477922 320058 477978
rect 350598 478294 350654 478350
rect 350722 478294 350778 478350
rect 350598 478170 350654 478226
rect 350722 478170 350778 478226
rect 350598 478046 350654 478102
rect 350722 478046 350778 478102
rect 350598 477922 350654 477978
rect 350722 477922 350778 477978
rect 381318 478294 381374 478350
rect 381442 478294 381498 478350
rect 381318 478170 381374 478226
rect 381442 478170 381498 478226
rect 381318 478046 381374 478102
rect 381442 478046 381498 478102
rect 381318 477922 381374 477978
rect 381442 477922 381498 477978
rect 412038 478294 412094 478350
rect 412162 478294 412218 478350
rect 412038 478170 412094 478226
rect 412162 478170 412218 478226
rect 412038 478046 412094 478102
rect 412162 478046 412218 478102
rect 412038 477922 412094 477978
rect 412162 477922 412218 477978
rect 442758 478294 442814 478350
rect 442882 478294 442938 478350
rect 442758 478170 442814 478226
rect 442882 478170 442938 478226
rect 442758 478046 442814 478102
rect 442882 478046 442938 478102
rect 442758 477922 442814 477978
rect 442882 477922 442938 477978
rect 303212 472562 303268 472618
rect 288204 431882 288260 431938
rect 285714 424294 285770 424350
rect 285838 424294 285894 424350
rect 285962 424294 286018 424350
rect 286086 424294 286142 424350
rect 285714 424170 285770 424226
rect 285838 424170 285894 424226
rect 285962 424170 286018 424226
rect 286086 424170 286142 424226
rect 285714 424046 285770 424102
rect 285838 424046 285894 424102
rect 285962 424046 286018 424102
rect 286086 424046 286142 424102
rect 285714 423922 285770 423978
rect 285838 423922 285894 423978
rect 285962 423922 286018 423978
rect 286086 423922 286142 423978
rect 285714 406294 285770 406350
rect 285838 406294 285894 406350
rect 285962 406294 286018 406350
rect 286086 406294 286142 406350
rect 285714 406170 285770 406226
rect 285838 406170 285894 406226
rect 285962 406170 286018 406226
rect 286086 406170 286142 406226
rect 285714 406046 285770 406102
rect 285838 406046 285894 406102
rect 285962 406046 286018 406102
rect 286086 406046 286142 406102
rect 285714 405922 285770 405978
rect 285838 405922 285894 405978
rect 285962 405922 286018 405978
rect 286086 405922 286142 405978
rect 285714 388294 285770 388350
rect 285838 388294 285894 388350
rect 285962 388294 286018 388350
rect 286086 388294 286142 388350
rect 285714 388170 285770 388226
rect 285838 388170 285894 388226
rect 285962 388170 286018 388226
rect 286086 388170 286142 388226
rect 285714 388046 285770 388102
rect 285838 388046 285894 388102
rect 285962 388046 286018 388102
rect 286086 388046 286142 388102
rect 285714 387922 285770 387978
rect 285838 387922 285894 387978
rect 285962 387922 286018 387978
rect 286086 387922 286142 387978
rect 285714 370294 285770 370350
rect 285838 370294 285894 370350
rect 285962 370294 286018 370350
rect 286086 370294 286142 370350
rect 285714 370170 285770 370226
rect 285838 370170 285894 370226
rect 285962 370170 286018 370226
rect 286086 370170 286142 370226
rect 285714 370046 285770 370102
rect 285838 370046 285894 370102
rect 285962 370046 286018 370102
rect 286086 370046 286142 370102
rect 285714 369922 285770 369978
rect 285838 369922 285894 369978
rect 285962 369922 286018 369978
rect 286086 369922 286142 369978
rect 285714 352294 285770 352350
rect 285838 352294 285894 352350
rect 285962 352294 286018 352350
rect 286086 352294 286142 352350
rect 285714 352170 285770 352226
rect 285838 352170 285894 352226
rect 285962 352170 286018 352226
rect 286086 352170 286142 352226
rect 285714 352046 285770 352102
rect 285838 352046 285894 352102
rect 285962 352046 286018 352102
rect 286086 352046 286142 352102
rect 285714 351922 285770 351978
rect 285838 351922 285894 351978
rect 285962 351922 286018 351978
rect 286086 351922 286142 351978
rect 284844 206342 284900 206398
rect 288092 339182 288148 339238
rect 285714 334294 285770 334350
rect 285838 334294 285894 334350
rect 285962 334294 286018 334350
rect 286086 334294 286142 334350
rect 285714 334170 285770 334226
rect 285838 334170 285894 334226
rect 285962 334170 286018 334226
rect 286086 334170 286142 334226
rect 285714 334046 285770 334102
rect 285838 334046 285894 334102
rect 285962 334046 286018 334102
rect 286086 334046 286142 334102
rect 285714 333922 285770 333978
rect 285838 333922 285894 333978
rect 285962 333922 286018 333978
rect 286086 333922 286142 333978
rect 285714 316294 285770 316350
rect 285838 316294 285894 316350
rect 285962 316294 286018 316350
rect 286086 316294 286142 316350
rect 285714 316170 285770 316226
rect 285838 316170 285894 316226
rect 285962 316170 286018 316226
rect 286086 316170 286142 316226
rect 285714 316046 285770 316102
rect 285838 316046 285894 316102
rect 285962 316046 286018 316102
rect 286086 316046 286142 316102
rect 285714 315922 285770 315978
rect 285838 315922 285894 315978
rect 285962 315922 286018 315978
rect 286086 315922 286142 315978
rect 285714 298294 285770 298350
rect 285838 298294 285894 298350
rect 285962 298294 286018 298350
rect 286086 298294 286142 298350
rect 285714 298170 285770 298226
rect 285838 298170 285894 298226
rect 285962 298170 286018 298226
rect 286086 298170 286142 298226
rect 285714 298046 285770 298102
rect 285838 298046 285894 298102
rect 285962 298046 286018 298102
rect 286086 298046 286142 298102
rect 285714 297922 285770 297978
rect 285838 297922 285894 297978
rect 285962 297922 286018 297978
rect 286086 297922 286142 297978
rect 285714 280294 285770 280350
rect 285838 280294 285894 280350
rect 285962 280294 286018 280350
rect 286086 280294 286142 280350
rect 285714 280170 285770 280226
rect 285838 280170 285894 280226
rect 285962 280170 286018 280226
rect 286086 280170 286142 280226
rect 285714 280046 285770 280102
rect 285838 280046 285894 280102
rect 285962 280046 286018 280102
rect 286086 280046 286142 280102
rect 285714 279922 285770 279978
rect 285838 279922 285894 279978
rect 285962 279922 286018 279978
rect 286086 279922 286142 279978
rect 285714 262294 285770 262350
rect 285838 262294 285894 262350
rect 285962 262294 286018 262350
rect 286086 262294 286142 262350
rect 285714 262170 285770 262226
rect 285838 262170 285894 262226
rect 285962 262170 286018 262226
rect 286086 262170 286142 262226
rect 285714 262046 285770 262102
rect 285838 262046 285894 262102
rect 285962 262046 286018 262102
rect 286086 262046 286142 262102
rect 285714 261922 285770 261978
rect 285838 261922 285894 261978
rect 285962 261922 286018 261978
rect 286086 261922 286142 261978
rect 285714 244294 285770 244350
rect 285838 244294 285894 244350
rect 285962 244294 286018 244350
rect 286086 244294 286142 244350
rect 285714 244170 285770 244226
rect 285838 244170 285894 244226
rect 285962 244170 286018 244226
rect 286086 244170 286142 244226
rect 285714 244046 285770 244102
rect 285838 244046 285894 244102
rect 285962 244046 286018 244102
rect 286086 244046 286142 244102
rect 285714 243922 285770 243978
rect 285838 243922 285894 243978
rect 285962 243922 286018 243978
rect 286086 243922 286142 243978
rect 285714 226294 285770 226350
rect 285838 226294 285894 226350
rect 285962 226294 286018 226350
rect 286086 226294 286142 226350
rect 285714 226170 285770 226226
rect 285838 226170 285894 226226
rect 285962 226170 286018 226226
rect 286086 226170 286142 226226
rect 285714 226046 285770 226102
rect 285838 226046 285894 226102
rect 285962 226046 286018 226102
rect 286086 226046 286142 226102
rect 285714 225922 285770 225978
rect 285838 225922 285894 225978
rect 285962 225922 286018 225978
rect 286086 225922 286142 225978
rect 285714 208294 285770 208350
rect 285838 208294 285894 208350
rect 285962 208294 286018 208350
rect 286086 208294 286142 208350
rect 285714 208170 285770 208226
rect 285838 208170 285894 208226
rect 285962 208170 286018 208226
rect 286086 208170 286142 208226
rect 285714 208046 285770 208102
rect 285838 208046 285894 208102
rect 285962 208046 286018 208102
rect 286086 208046 286142 208102
rect 285714 207922 285770 207978
rect 285838 207922 285894 207978
rect 285962 207922 286018 207978
rect 286086 207922 286142 207978
rect 285714 190294 285770 190350
rect 285838 190294 285894 190350
rect 285962 190294 286018 190350
rect 286086 190294 286142 190350
rect 285714 190170 285770 190226
rect 285838 190170 285894 190226
rect 285962 190170 286018 190226
rect 286086 190170 286142 190226
rect 285714 190046 285770 190102
rect 285838 190046 285894 190102
rect 285962 190046 286018 190102
rect 286086 190046 286142 190102
rect 285714 189922 285770 189978
rect 285838 189922 285894 189978
rect 285962 189922 286018 189978
rect 286086 189922 286142 189978
rect 285714 172294 285770 172350
rect 285838 172294 285894 172350
rect 285962 172294 286018 172350
rect 286086 172294 286142 172350
rect 285714 172170 285770 172226
rect 285838 172170 285894 172226
rect 285962 172170 286018 172226
rect 286086 172170 286142 172226
rect 285714 172046 285770 172102
rect 285838 172046 285894 172102
rect 285962 172046 286018 172102
rect 286086 172046 286142 172102
rect 285714 171922 285770 171978
rect 285838 171922 285894 171978
rect 285962 171922 286018 171978
rect 286086 171922 286142 171978
rect 285714 154294 285770 154350
rect 285838 154294 285894 154350
rect 285962 154294 286018 154350
rect 286086 154294 286142 154350
rect 285714 154170 285770 154226
rect 285838 154170 285894 154226
rect 285962 154170 286018 154226
rect 286086 154170 286142 154226
rect 285714 154046 285770 154102
rect 285838 154046 285894 154102
rect 285962 154046 286018 154102
rect 286086 154046 286142 154102
rect 285714 153922 285770 153978
rect 285838 153922 285894 153978
rect 285962 153922 286018 153978
rect 286086 153922 286142 153978
rect 285714 136294 285770 136350
rect 285838 136294 285894 136350
rect 285962 136294 286018 136350
rect 286086 136294 286142 136350
rect 285714 136170 285770 136226
rect 285838 136170 285894 136226
rect 285962 136170 286018 136226
rect 286086 136170 286142 136226
rect 285714 136046 285770 136102
rect 285838 136046 285894 136102
rect 285962 136046 286018 136102
rect 286086 136046 286142 136102
rect 285714 135922 285770 135978
rect 285838 135922 285894 135978
rect 285962 135922 286018 135978
rect 286086 135922 286142 135978
rect 285714 118294 285770 118350
rect 285838 118294 285894 118350
rect 285962 118294 286018 118350
rect 286086 118294 286142 118350
rect 285714 118170 285770 118226
rect 285838 118170 285894 118226
rect 285962 118170 286018 118226
rect 286086 118170 286142 118226
rect 285714 118046 285770 118102
rect 285838 118046 285894 118102
rect 285962 118046 286018 118102
rect 286086 118046 286142 118102
rect 285714 117922 285770 117978
rect 285838 117922 285894 117978
rect 285962 117922 286018 117978
rect 286086 117922 286142 117978
rect 285714 100294 285770 100350
rect 285838 100294 285894 100350
rect 285962 100294 286018 100350
rect 286086 100294 286142 100350
rect 285714 100170 285770 100226
rect 285838 100170 285894 100226
rect 285962 100170 286018 100226
rect 286086 100170 286142 100226
rect 285714 100046 285770 100102
rect 285838 100046 285894 100102
rect 285962 100046 286018 100102
rect 286086 100046 286142 100102
rect 285714 99922 285770 99978
rect 285838 99922 285894 99978
rect 285962 99922 286018 99978
rect 286086 99922 286142 99978
rect 285714 82294 285770 82350
rect 285838 82294 285894 82350
rect 285962 82294 286018 82350
rect 286086 82294 286142 82350
rect 285714 82170 285770 82226
rect 285838 82170 285894 82226
rect 285962 82170 286018 82226
rect 286086 82170 286142 82226
rect 285714 82046 285770 82102
rect 285838 82046 285894 82102
rect 285962 82046 286018 82102
rect 286086 82046 286142 82102
rect 285714 81922 285770 81978
rect 285838 81922 285894 81978
rect 285962 81922 286018 81978
rect 286086 81922 286142 81978
rect 285714 64294 285770 64350
rect 285838 64294 285894 64350
rect 285962 64294 286018 64350
rect 286086 64294 286142 64350
rect 285714 64170 285770 64226
rect 285838 64170 285894 64226
rect 285962 64170 286018 64226
rect 286086 64170 286142 64226
rect 285714 64046 285770 64102
rect 285838 64046 285894 64102
rect 285962 64046 286018 64102
rect 286086 64046 286142 64102
rect 285714 63922 285770 63978
rect 285838 63922 285894 63978
rect 285962 63922 286018 63978
rect 286086 63922 286142 63978
rect 285714 46294 285770 46350
rect 285838 46294 285894 46350
rect 285962 46294 286018 46350
rect 286086 46294 286142 46350
rect 285714 46170 285770 46226
rect 285838 46170 285894 46226
rect 285962 46170 286018 46226
rect 286086 46170 286142 46226
rect 285714 46046 285770 46102
rect 285838 46046 285894 46102
rect 285962 46046 286018 46102
rect 286086 46046 286142 46102
rect 285714 45922 285770 45978
rect 285838 45922 285894 45978
rect 285962 45922 286018 45978
rect 286086 45922 286142 45978
rect 285714 28294 285770 28350
rect 285838 28294 285894 28350
rect 285962 28294 286018 28350
rect 286086 28294 286142 28350
rect 285714 28170 285770 28226
rect 285838 28170 285894 28226
rect 285962 28170 286018 28226
rect 286086 28170 286142 28226
rect 285714 28046 285770 28102
rect 285838 28046 285894 28102
rect 285962 28046 286018 28102
rect 286086 28046 286142 28102
rect 285714 27922 285770 27978
rect 285838 27922 285894 27978
rect 285962 27922 286018 27978
rect 286086 27922 286142 27978
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 285714 10294 285770 10350
rect 285838 10294 285894 10350
rect 285962 10294 286018 10350
rect 286086 10294 286142 10350
rect 285714 10170 285770 10226
rect 285838 10170 285894 10226
rect 285962 10170 286018 10226
rect 286086 10170 286142 10226
rect 285714 10046 285770 10102
rect 285838 10046 285894 10102
rect 285962 10046 286018 10102
rect 286086 10046 286142 10102
rect 285714 9922 285770 9978
rect 285838 9922 285894 9978
rect 285962 9922 286018 9978
rect 286086 9922 286142 9978
rect 289772 427022 289828 427078
rect 289884 377882 289940 377938
rect 289772 345482 289828 345538
rect 288316 326042 288372 326098
rect 289884 317762 289940 317818
rect 296604 430802 296660 430858
rect 293132 377702 293188 377758
rect 291564 285182 291620 285238
rect 294812 425402 294868 425458
rect 295260 373742 295316 373798
rect 295036 368702 295092 368758
rect 294924 360242 294980 360298
rect 294812 348542 294868 348598
rect 298172 430082 298228 430138
rect 298060 426842 298116 426898
rect 296604 377522 296660 377578
rect 296492 345122 296548 345178
rect 293244 332522 293300 332578
rect 293244 314162 293300 314218
rect 299964 430982 300020 431038
rect 298396 402722 298452 402778
rect 298508 428462 298564 428518
rect 298620 404522 298676 404578
rect 299852 425042 299908 425098
rect 298732 398042 298788 398098
rect 298284 337382 298340 337438
rect 299852 332342 299908 332398
rect 300860 427382 300916 427438
rect 301532 427382 301588 427438
rect 300972 425222 301028 425278
rect 304518 472294 304574 472350
rect 304642 472294 304698 472350
rect 304518 472170 304574 472226
rect 304642 472170 304698 472226
rect 304518 472046 304574 472102
rect 304642 472046 304698 472102
rect 304518 471922 304574 471978
rect 304642 471922 304698 471978
rect 335238 472294 335294 472350
rect 335362 472294 335418 472350
rect 335238 472170 335294 472226
rect 335362 472170 335418 472226
rect 335238 472046 335294 472102
rect 335362 472046 335418 472102
rect 335238 471922 335294 471978
rect 335362 471922 335418 471978
rect 365958 472294 366014 472350
rect 366082 472294 366138 472350
rect 365958 472170 366014 472226
rect 366082 472170 366138 472226
rect 365958 472046 366014 472102
rect 366082 472046 366138 472102
rect 365958 471922 366014 471978
rect 366082 471922 366138 471978
rect 396678 472294 396734 472350
rect 396802 472294 396858 472350
rect 396678 472170 396734 472226
rect 396802 472170 396858 472226
rect 396678 472046 396734 472102
rect 396802 472046 396858 472102
rect 396678 471922 396734 471978
rect 396802 471922 396858 471978
rect 427398 472294 427454 472350
rect 427522 472294 427578 472350
rect 427398 472170 427454 472226
rect 427522 472170 427578 472226
rect 427398 472046 427454 472102
rect 427522 472046 427578 472102
rect 427398 471922 427454 471978
rect 427522 471922 427578 471978
rect 319878 460294 319934 460350
rect 320002 460294 320058 460350
rect 319878 460170 319934 460226
rect 320002 460170 320058 460226
rect 319878 460046 319934 460102
rect 320002 460046 320058 460102
rect 319878 459922 319934 459978
rect 320002 459922 320058 459978
rect 350598 460294 350654 460350
rect 350722 460294 350778 460350
rect 350598 460170 350654 460226
rect 350722 460170 350778 460226
rect 350598 460046 350654 460102
rect 350722 460046 350778 460102
rect 350598 459922 350654 459978
rect 350722 459922 350778 459978
rect 381318 460294 381374 460350
rect 381442 460294 381498 460350
rect 381318 460170 381374 460226
rect 381442 460170 381498 460226
rect 381318 460046 381374 460102
rect 381442 460046 381498 460102
rect 381318 459922 381374 459978
rect 381442 459922 381498 459978
rect 412038 460294 412094 460350
rect 412162 460294 412218 460350
rect 412038 460170 412094 460226
rect 412162 460170 412218 460226
rect 412038 460046 412094 460102
rect 412162 460046 412218 460102
rect 412038 459922 412094 459978
rect 412162 459922 412218 459978
rect 442758 460294 442814 460350
rect 442882 460294 442938 460350
rect 442758 460170 442814 460226
rect 442882 460170 442938 460226
rect 442758 460046 442814 460102
rect 442882 460046 442938 460102
rect 442758 459922 442814 459978
rect 442882 459922 442938 459978
rect 304518 454294 304574 454350
rect 304642 454294 304698 454350
rect 304518 454170 304574 454226
rect 304642 454170 304698 454226
rect 304518 454046 304574 454102
rect 304642 454046 304698 454102
rect 304518 453922 304574 453978
rect 304642 453922 304698 453978
rect 335238 454294 335294 454350
rect 335362 454294 335418 454350
rect 335238 454170 335294 454226
rect 335362 454170 335418 454226
rect 335238 454046 335294 454102
rect 335362 454046 335418 454102
rect 335238 453922 335294 453978
rect 335362 453922 335418 453978
rect 365958 454294 366014 454350
rect 366082 454294 366138 454350
rect 365958 454170 366014 454226
rect 366082 454170 366138 454226
rect 365958 454046 366014 454102
rect 366082 454046 366138 454102
rect 365958 453922 366014 453978
rect 366082 453922 366138 453978
rect 396678 454294 396734 454350
rect 396802 454294 396858 454350
rect 396678 454170 396734 454226
rect 396802 454170 396858 454226
rect 396678 454046 396734 454102
rect 396802 454046 396858 454102
rect 396678 453922 396734 453978
rect 396802 453922 396858 453978
rect 427398 454294 427454 454350
rect 427522 454294 427578 454350
rect 427398 454170 427454 454226
rect 427522 454170 427578 454226
rect 427398 454046 427454 454102
rect 427522 454046 427578 454102
rect 427398 453922 427454 453978
rect 427522 453922 427578 453978
rect 319878 442294 319934 442350
rect 320002 442294 320058 442350
rect 319878 442170 319934 442226
rect 320002 442170 320058 442226
rect 319878 442046 319934 442102
rect 320002 442046 320058 442102
rect 319878 441922 319934 441978
rect 320002 441922 320058 441978
rect 350598 442294 350654 442350
rect 350722 442294 350778 442350
rect 350598 442170 350654 442226
rect 350722 442170 350778 442226
rect 350598 442046 350654 442102
rect 350722 442046 350778 442102
rect 350598 441922 350654 441978
rect 350722 441922 350778 441978
rect 381318 442294 381374 442350
rect 381442 442294 381498 442350
rect 381318 442170 381374 442226
rect 381442 442170 381498 442226
rect 381318 442046 381374 442102
rect 381442 442046 381498 442102
rect 381318 441922 381374 441978
rect 381442 441922 381498 441978
rect 412038 442294 412094 442350
rect 412162 442294 412218 442350
rect 412038 442170 412094 442226
rect 412162 442170 412218 442226
rect 412038 442046 412094 442102
rect 412162 442046 412218 442102
rect 412038 441922 412094 441978
rect 412162 441922 412218 441978
rect 442758 442294 442814 442350
rect 442882 442294 442938 442350
rect 442758 442170 442814 442226
rect 442882 442170 442938 442226
rect 442758 442046 442814 442102
rect 442882 442046 442938 442102
rect 442758 441922 442814 441978
rect 442882 441922 442938 441978
rect 304518 436294 304574 436350
rect 304642 436294 304698 436350
rect 304518 436170 304574 436226
rect 304642 436170 304698 436226
rect 304518 436046 304574 436102
rect 304642 436046 304698 436102
rect 304518 435922 304574 435978
rect 304642 435922 304698 435978
rect 335238 436294 335294 436350
rect 335362 436294 335418 436350
rect 335238 436170 335294 436226
rect 335362 436170 335418 436226
rect 335238 436046 335294 436102
rect 335362 436046 335418 436102
rect 335238 435922 335294 435978
rect 335362 435922 335418 435978
rect 365958 436294 366014 436350
rect 366082 436294 366138 436350
rect 365958 436170 366014 436226
rect 366082 436170 366138 436226
rect 365958 436046 366014 436102
rect 366082 436046 366138 436102
rect 365958 435922 366014 435978
rect 366082 435922 366138 435978
rect 396678 436294 396734 436350
rect 396802 436294 396858 436350
rect 396678 436170 396734 436226
rect 396802 436170 396858 436226
rect 396678 436046 396734 436102
rect 396802 436046 396858 436102
rect 396678 435922 396734 435978
rect 396802 435922 396858 435978
rect 427398 436294 427454 436350
rect 427522 436294 427578 436350
rect 427398 436170 427454 436226
rect 427522 436170 427578 436226
rect 427398 436046 427454 436102
rect 427522 436046 427578 436102
rect 427398 435922 427454 435978
rect 427522 435922 427578 435978
rect 452732 433322 452788 433378
rect 457772 548162 457828 548218
rect 319878 424294 319934 424350
rect 320002 424294 320058 424350
rect 319878 424170 319934 424226
rect 320002 424170 320058 424226
rect 319878 424046 319934 424102
rect 320002 424046 320058 424102
rect 319878 423922 319934 423978
rect 320002 423922 320058 423978
rect 350598 424294 350654 424350
rect 350722 424294 350778 424350
rect 350598 424170 350654 424226
rect 350722 424170 350778 424226
rect 350598 424046 350654 424102
rect 350722 424046 350778 424102
rect 350598 423922 350654 423978
rect 350722 423922 350778 423978
rect 381318 424294 381374 424350
rect 381442 424294 381498 424350
rect 381318 424170 381374 424226
rect 381442 424170 381498 424226
rect 381318 424046 381374 424102
rect 381442 424046 381498 424102
rect 381318 423922 381374 423978
rect 381442 423922 381498 423978
rect 412038 424294 412094 424350
rect 412162 424294 412218 424350
rect 412038 424170 412094 424226
rect 412162 424170 412218 424226
rect 412038 424046 412094 424102
rect 412162 424046 412218 424102
rect 412038 423922 412094 423978
rect 412162 423922 412218 423978
rect 442758 424294 442814 424350
rect 442882 424294 442938 424350
rect 442758 424170 442814 424226
rect 442882 424170 442938 424226
rect 442758 424046 442814 424102
rect 442882 424046 442938 424102
rect 442758 423922 442814 423978
rect 442882 423922 442938 423978
rect 304518 418294 304574 418350
rect 304642 418294 304698 418350
rect 304518 418170 304574 418226
rect 304642 418170 304698 418226
rect 304518 418046 304574 418102
rect 304642 418046 304698 418102
rect 304518 417922 304574 417978
rect 304642 417922 304698 417978
rect 335238 418294 335294 418350
rect 335362 418294 335418 418350
rect 335238 418170 335294 418226
rect 335362 418170 335418 418226
rect 335238 418046 335294 418102
rect 335362 418046 335418 418102
rect 335238 417922 335294 417978
rect 335362 417922 335418 417978
rect 365958 418294 366014 418350
rect 366082 418294 366138 418350
rect 365958 418170 366014 418226
rect 366082 418170 366138 418226
rect 365958 418046 366014 418102
rect 366082 418046 366138 418102
rect 365958 417922 366014 417978
rect 366082 417922 366138 417978
rect 396678 418294 396734 418350
rect 396802 418294 396858 418350
rect 396678 418170 396734 418226
rect 396802 418170 396858 418226
rect 396678 418046 396734 418102
rect 396802 418046 396858 418102
rect 396678 417922 396734 417978
rect 396802 417922 396858 417978
rect 427398 418294 427454 418350
rect 427522 418294 427578 418350
rect 427398 418170 427454 418226
rect 427522 418170 427578 418226
rect 427398 418046 427454 418102
rect 427522 418046 427578 418102
rect 427398 417922 427454 417978
rect 427522 417922 427578 417978
rect 319878 406294 319934 406350
rect 320002 406294 320058 406350
rect 319878 406170 319934 406226
rect 320002 406170 320058 406226
rect 319878 406046 319934 406102
rect 320002 406046 320058 406102
rect 319878 405922 319934 405978
rect 320002 405922 320058 405978
rect 350598 406294 350654 406350
rect 350722 406294 350778 406350
rect 350598 406170 350654 406226
rect 350722 406170 350778 406226
rect 350598 406046 350654 406102
rect 350722 406046 350778 406102
rect 350598 405922 350654 405978
rect 350722 405922 350778 405978
rect 381318 406294 381374 406350
rect 381442 406294 381498 406350
rect 381318 406170 381374 406226
rect 381442 406170 381498 406226
rect 381318 406046 381374 406102
rect 381442 406046 381498 406102
rect 381318 405922 381374 405978
rect 381442 405922 381498 405978
rect 412038 406294 412094 406350
rect 412162 406294 412218 406350
rect 412038 406170 412094 406226
rect 412162 406170 412218 406226
rect 412038 406046 412094 406102
rect 412162 406046 412218 406102
rect 412038 405922 412094 405978
rect 412162 405922 412218 405978
rect 442758 406294 442814 406350
rect 442882 406294 442938 406350
rect 442758 406170 442814 406226
rect 442882 406170 442938 406226
rect 442758 406046 442814 406102
rect 442882 406046 442938 406102
rect 442758 405922 442814 405978
rect 442882 405922 442938 405978
rect 303212 404342 303268 404398
rect 312714 400294 312770 400350
rect 312838 400294 312894 400350
rect 312962 400294 313018 400350
rect 313086 400294 313142 400350
rect 312714 400170 312770 400226
rect 312838 400170 312894 400226
rect 312962 400170 313018 400226
rect 313086 400170 313142 400226
rect 312714 400046 312770 400102
rect 312838 400046 312894 400102
rect 312962 400046 313018 400102
rect 313086 400046 313142 400102
rect 312714 399922 312770 399978
rect 312838 399922 312894 399978
rect 312962 399922 313018 399978
rect 313086 399922 313142 399978
rect 312714 382294 312770 382350
rect 312838 382294 312894 382350
rect 312962 382294 313018 382350
rect 313086 382294 313142 382350
rect 312714 382170 312770 382226
rect 312838 382170 312894 382226
rect 312962 382170 313018 382226
rect 313086 382170 313142 382226
rect 312714 382046 312770 382102
rect 312838 382046 312894 382102
rect 312962 382046 313018 382102
rect 313086 382046 313142 382102
rect 312714 381922 312770 381978
rect 312838 381922 312894 381978
rect 312962 381922 313018 381978
rect 313086 381922 313142 381978
rect 301932 370294 301988 370350
rect 302056 370294 302112 370350
rect 302180 370294 302236 370350
rect 302304 370294 302360 370350
rect 301932 370170 301988 370226
rect 302056 370170 302112 370226
rect 302180 370170 302236 370226
rect 302304 370170 302360 370226
rect 301932 370046 301988 370102
rect 302056 370046 302112 370102
rect 302180 370046 302236 370102
rect 302304 370046 302360 370102
rect 301932 369922 301988 369978
rect 302056 369922 302112 369978
rect 302180 369922 302236 369978
rect 302304 369922 302360 369978
rect 302732 364294 302788 364350
rect 302856 364294 302912 364350
rect 302980 364294 303036 364350
rect 303104 364294 303160 364350
rect 302732 364170 302788 364226
rect 302856 364170 302912 364226
rect 302980 364170 303036 364226
rect 303104 364170 303160 364226
rect 302732 364046 302788 364102
rect 302856 364046 302912 364102
rect 302980 364046 303036 364102
rect 303104 364046 303160 364102
rect 302732 363922 302788 363978
rect 302856 363922 302912 363978
rect 302980 363922 303036 363978
rect 303104 363922 303160 363978
rect 312714 364294 312770 364350
rect 312838 364294 312894 364350
rect 312962 364294 313018 364350
rect 313086 364294 313142 364350
rect 312714 364170 312770 364226
rect 312838 364170 312894 364226
rect 312962 364170 313018 364226
rect 313086 364170 313142 364226
rect 312714 364046 312770 364102
rect 312838 364046 312894 364102
rect 312962 364046 313018 364102
rect 313086 364046 313142 364102
rect 312714 363922 312770 363978
rect 312838 363922 312894 363978
rect 312962 363922 313018 363978
rect 313086 363922 313142 363978
rect 301932 352294 301988 352350
rect 302056 352294 302112 352350
rect 302180 352294 302236 352350
rect 302304 352294 302360 352350
rect 301932 352170 301988 352226
rect 302056 352170 302112 352226
rect 302180 352170 302236 352226
rect 302304 352170 302360 352226
rect 301932 352046 301988 352102
rect 302056 352046 302112 352102
rect 302180 352046 302236 352102
rect 302304 352046 302360 352102
rect 301932 351922 301988 351978
rect 302056 351922 302112 351978
rect 302180 351922 302236 351978
rect 302304 351922 302360 351978
rect 302732 346294 302788 346350
rect 302856 346294 302912 346350
rect 302980 346294 303036 346350
rect 303104 346294 303160 346350
rect 302732 346170 302788 346226
rect 302856 346170 302912 346226
rect 302980 346170 303036 346226
rect 303104 346170 303160 346226
rect 302732 346046 302788 346102
rect 302856 346046 302912 346102
rect 302980 346046 303036 346102
rect 303104 346046 303160 346102
rect 302732 345922 302788 345978
rect 302856 345922 302912 345978
rect 302980 345922 303036 345978
rect 303104 345922 303160 345978
rect 312714 346294 312770 346350
rect 312838 346294 312894 346350
rect 312962 346294 313018 346350
rect 313086 346294 313142 346350
rect 312714 346170 312770 346226
rect 312838 346170 312894 346226
rect 312962 346170 313018 346226
rect 313086 346170 313142 346226
rect 312714 346046 312770 346102
rect 312838 346046 312894 346102
rect 312962 346046 313018 346102
rect 313086 346046 313142 346102
rect 312714 345922 312770 345978
rect 312838 345922 312894 345978
rect 312962 345922 313018 345978
rect 313086 345922 313142 345978
rect 301084 340262 301140 340318
rect 300860 340082 300916 340138
rect 301932 334294 301988 334350
rect 302056 334294 302112 334350
rect 302180 334294 302236 334350
rect 302304 334294 302360 334350
rect 301932 334170 301988 334226
rect 302056 334170 302112 334226
rect 302180 334170 302236 334226
rect 302304 334170 302360 334226
rect 301932 334046 301988 334102
rect 302056 334046 302112 334102
rect 302180 334046 302236 334102
rect 302304 334046 302360 334102
rect 301932 333922 301988 333978
rect 302056 333922 302112 333978
rect 302180 333922 302236 333978
rect 302304 333922 302360 333978
rect 302732 328294 302788 328350
rect 302856 328294 302912 328350
rect 302980 328294 303036 328350
rect 303104 328294 303160 328350
rect 302732 328170 302788 328226
rect 302856 328170 302912 328226
rect 302980 328170 303036 328226
rect 303104 328170 303160 328226
rect 302732 328046 302788 328102
rect 302856 328046 302912 328102
rect 302980 328046 303036 328102
rect 303104 328046 303160 328102
rect 302732 327922 302788 327978
rect 302856 327922 302912 327978
rect 302980 327922 303036 327978
rect 303104 327922 303160 327978
rect 312714 328294 312770 328350
rect 312838 328294 312894 328350
rect 312962 328294 313018 328350
rect 313086 328294 313142 328350
rect 312714 328170 312770 328226
rect 312838 328170 312894 328226
rect 312962 328170 313018 328226
rect 313086 328170 313142 328226
rect 312714 328046 312770 328102
rect 312838 328046 312894 328102
rect 312962 328046 313018 328102
rect 313086 328046 313142 328102
rect 312714 327922 312770 327978
rect 312838 327922 312894 327978
rect 312962 327922 313018 327978
rect 313086 327922 313142 327978
rect 301932 316294 301988 316350
rect 302056 316294 302112 316350
rect 302180 316294 302236 316350
rect 302304 316294 302360 316350
rect 301932 316170 301988 316226
rect 302056 316170 302112 316226
rect 302180 316170 302236 316226
rect 302304 316170 302360 316226
rect 301932 316046 301988 316102
rect 302056 316046 302112 316102
rect 302180 316046 302236 316102
rect 302304 316046 302360 316102
rect 301932 315922 301988 315978
rect 302056 315922 302112 315978
rect 302180 315922 302236 315978
rect 302304 315922 302360 315978
rect 302732 310294 302788 310350
rect 302856 310294 302912 310350
rect 302980 310294 303036 310350
rect 303104 310294 303160 310350
rect 302732 310170 302788 310226
rect 302856 310170 302912 310226
rect 302980 310170 303036 310226
rect 303104 310170 303160 310226
rect 302732 310046 302788 310102
rect 302856 310046 302912 310102
rect 302980 310046 303036 310102
rect 303104 310046 303160 310102
rect 302732 309922 302788 309978
rect 302856 309922 302912 309978
rect 302980 309922 303036 309978
rect 303104 309922 303160 309978
rect 312714 310294 312770 310350
rect 312838 310294 312894 310350
rect 312962 310294 313018 310350
rect 313086 310294 313142 310350
rect 312714 310170 312770 310226
rect 312838 310170 312894 310226
rect 312962 310170 313018 310226
rect 313086 310170 313142 310226
rect 312714 310046 312770 310102
rect 312838 310046 312894 310102
rect 312962 310046 313018 310102
rect 313086 310046 313142 310102
rect 312714 309922 312770 309978
rect 312838 309922 312894 309978
rect 312962 309922 313018 309978
rect 313086 309922 313142 309978
rect 301932 298294 301988 298350
rect 302056 298294 302112 298350
rect 302180 298294 302236 298350
rect 302304 298294 302360 298350
rect 301932 298170 301988 298226
rect 302056 298170 302112 298226
rect 302180 298170 302236 298226
rect 302304 298170 302360 298226
rect 301932 298046 301988 298102
rect 302056 298046 302112 298102
rect 302180 298046 302236 298102
rect 302304 298046 302360 298102
rect 301932 297922 301988 297978
rect 302056 297922 302112 297978
rect 302180 297922 302236 297978
rect 302304 297922 302360 297978
rect 302732 292294 302788 292350
rect 302856 292294 302912 292350
rect 302980 292294 303036 292350
rect 303104 292294 303160 292350
rect 302732 292170 302788 292226
rect 302856 292170 302912 292226
rect 302980 292170 303036 292226
rect 303104 292170 303160 292226
rect 302732 292046 302788 292102
rect 302856 292046 302912 292102
rect 302980 292046 303036 292102
rect 303104 292046 303160 292102
rect 302732 291922 302788 291978
rect 302856 291922 302912 291978
rect 302980 291922 303036 291978
rect 303104 291922 303160 291978
rect 312714 292294 312770 292350
rect 312838 292294 312894 292350
rect 312962 292294 313018 292350
rect 313086 292294 313142 292350
rect 312714 292170 312770 292226
rect 312838 292170 312894 292226
rect 312962 292170 313018 292226
rect 313086 292170 313142 292226
rect 312714 292046 312770 292102
rect 312838 292046 312894 292102
rect 312962 292046 313018 292102
rect 313086 292046 313142 292102
rect 312714 291922 312770 291978
rect 312838 291922 312894 291978
rect 312962 291922 313018 291978
rect 313086 291922 313142 291978
rect 304780 142082 304836 142138
rect 303996 140822 304052 140878
rect 299964 127502 300020 127558
rect 312714 274294 312770 274350
rect 312838 274294 312894 274350
rect 312962 274294 313018 274350
rect 313086 274294 313142 274350
rect 312714 274170 312770 274226
rect 312838 274170 312894 274226
rect 312962 274170 313018 274226
rect 313086 274170 313142 274226
rect 312714 274046 312770 274102
rect 312838 274046 312894 274102
rect 312962 274046 313018 274102
rect 313086 274046 313142 274102
rect 312714 273922 312770 273978
rect 312838 273922 312894 273978
rect 312962 273922 313018 273978
rect 313086 273922 313142 273978
rect 312714 256294 312770 256350
rect 312838 256294 312894 256350
rect 312962 256294 313018 256350
rect 313086 256294 313142 256350
rect 312714 256170 312770 256226
rect 312838 256170 312894 256226
rect 312962 256170 313018 256226
rect 313086 256170 313142 256226
rect 312714 256046 312770 256102
rect 312838 256046 312894 256102
rect 312962 256046 313018 256102
rect 313086 256046 313142 256102
rect 312714 255922 312770 255978
rect 312838 255922 312894 255978
rect 312962 255922 313018 255978
rect 313086 255922 313142 255978
rect 312714 238294 312770 238350
rect 312838 238294 312894 238350
rect 312962 238294 313018 238350
rect 313086 238294 313142 238350
rect 312714 238170 312770 238226
rect 312838 238170 312894 238226
rect 312962 238170 313018 238226
rect 313086 238170 313142 238226
rect 312714 238046 312770 238102
rect 312838 238046 312894 238102
rect 312962 238046 313018 238102
rect 313086 238046 313142 238102
rect 312714 237922 312770 237978
rect 312838 237922 312894 237978
rect 312962 237922 313018 237978
rect 313086 237922 313142 237978
rect 312714 220294 312770 220350
rect 312838 220294 312894 220350
rect 312962 220294 313018 220350
rect 313086 220294 313142 220350
rect 312714 220170 312770 220226
rect 312838 220170 312894 220226
rect 312962 220170 313018 220226
rect 313086 220170 313142 220226
rect 312714 220046 312770 220102
rect 312838 220046 312894 220102
rect 312962 220046 313018 220102
rect 313086 220046 313142 220102
rect 312714 219922 312770 219978
rect 312838 219922 312894 219978
rect 312962 219922 313018 219978
rect 313086 219922 313142 219978
rect 312714 202294 312770 202350
rect 312838 202294 312894 202350
rect 312962 202294 313018 202350
rect 313086 202294 313142 202350
rect 312714 202170 312770 202226
rect 312838 202170 312894 202226
rect 312962 202170 313018 202226
rect 313086 202170 313142 202226
rect 312714 202046 312770 202102
rect 312838 202046 312894 202102
rect 312962 202046 313018 202102
rect 313086 202046 313142 202102
rect 312714 201922 312770 201978
rect 312838 201922 312894 201978
rect 312962 201922 313018 201978
rect 313086 201922 313142 201978
rect 312714 184294 312770 184350
rect 312838 184294 312894 184350
rect 312962 184294 313018 184350
rect 313086 184294 313142 184350
rect 312714 184170 312770 184226
rect 312838 184170 312894 184226
rect 312962 184170 313018 184226
rect 313086 184170 313142 184226
rect 312714 184046 312770 184102
rect 312838 184046 312894 184102
rect 312962 184046 313018 184102
rect 313086 184046 313142 184102
rect 312714 183922 312770 183978
rect 312838 183922 312894 183978
rect 312962 183922 313018 183978
rect 313086 183922 313142 183978
rect 312714 166294 312770 166350
rect 312838 166294 312894 166350
rect 312962 166294 313018 166350
rect 313086 166294 313142 166350
rect 312714 166170 312770 166226
rect 312838 166170 312894 166226
rect 312962 166170 313018 166226
rect 313086 166170 313142 166226
rect 312714 166046 312770 166102
rect 312838 166046 312894 166102
rect 312962 166046 313018 166102
rect 313086 166046 313142 166102
rect 312714 165922 312770 165978
rect 312838 165922 312894 165978
rect 312962 165922 313018 165978
rect 313086 165922 313142 165978
rect 312714 148294 312770 148350
rect 312838 148294 312894 148350
rect 312962 148294 313018 148350
rect 313086 148294 313142 148350
rect 312714 148170 312770 148226
rect 312838 148170 312894 148226
rect 312962 148170 313018 148226
rect 313086 148170 313142 148226
rect 312714 148046 312770 148102
rect 312838 148046 312894 148102
rect 312962 148046 313018 148102
rect 313086 148046 313142 148102
rect 312714 147922 312770 147978
rect 312838 147922 312894 147978
rect 312962 147922 313018 147978
rect 313086 147922 313142 147978
rect 316434 388294 316490 388350
rect 316558 388294 316614 388350
rect 316682 388294 316738 388350
rect 316806 388294 316862 388350
rect 316434 388170 316490 388226
rect 316558 388170 316614 388226
rect 316682 388170 316738 388226
rect 316806 388170 316862 388226
rect 316434 388046 316490 388102
rect 316558 388046 316614 388102
rect 316682 388046 316738 388102
rect 316806 388046 316862 388102
rect 316434 387922 316490 387978
rect 316558 387922 316614 387978
rect 316682 387922 316738 387978
rect 316806 387922 316862 387978
rect 316434 370294 316490 370350
rect 316558 370294 316614 370350
rect 316682 370294 316738 370350
rect 316806 370294 316862 370350
rect 316434 370170 316490 370226
rect 316558 370170 316614 370226
rect 316682 370170 316738 370226
rect 316806 370170 316862 370226
rect 316434 370046 316490 370102
rect 316558 370046 316614 370102
rect 316682 370046 316738 370102
rect 316806 370046 316862 370102
rect 316434 369922 316490 369978
rect 316558 369922 316614 369978
rect 316682 369922 316738 369978
rect 316806 369922 316862 369978
rect 316434 352294 316490 352350
rect 316558 352294 316614 352350
rect 316682 352294 316738 352350
rect 316806 352294 316862 352350
rect 316434 352170 316490 352226
rect 316558 352170 316614 352226
rect 316682 352170 316738 352226
rect 316806 352170 316862 352226
rect 316434 352046 316490 352102
rect 316558 352046 316614 352102
rect 316682 352046 316738 352102
rect 316806 352046 316862 352102
rect 316434 351922 316490 351978
rect 316558 351922 316614 351978
rect 316682 351922 316738 351978
rect 316806 351922 316862 351978
rect 316434 334294 316490 334350
rect 316558 334294 316614 334350
rect 316682 334294 316738 334350
rect 316806 334294 316862 334350
rect 316434 334170 316490 334226
rect 316558 334170 316614 334226
rect 316682 334170 316738 334226
rect 316806 334170 316862 334226
rect 316434 334046 316490 334102
rect 316558 334046 316614 334102
rect 316682 334046 316738 334102
rect 316806 334046 316862 334102
rect 316434 333922 316490 333978
rect 316558 333922 316614 333978
rect 316682 333922 316738 333978
rect 316806 333922 316862 333978
rect 316434 316294 316490 316350
rect 316558 316294 316614 316350
rect 316682 316294 316738 316350
rect 316806 316294 316862 316350
rect 316434 316170 316490 316226
rect 316558 316170 316614 316226
rect 316682 316170 316738 316226
rect 316806 316170 316862 316226
rect 316434 316046 316490 316102
rect 316558 316046 316614 316102
rect 316682 316046 316738 316102
rect 316806 316046 316862 316102
rect 316434 315922 316490 315978
rect 316558 315922 316614 315978
rect 316682 315922 316738 315978
rect 316806 315922 316862 315978
rect 316434 298294 316490 298350
rect 316558 298294 316614 298350
rect 316682 298294 316738 298350
rect 316806 298294 316862 298350
rect 316434 298170 316490 298226
rect 316558 298170 316614 298226
rect 316682 298170 316738 298226
rect 316806 298170 316862 298226
rect 316434 298046 316490 298102
rect 316558 298046 316614 298102
rect 316682 298046 316738 298102
rect 316806 298046 316862 298102
rect 316434 297922 316490 297978
rect 316558 297922 316614 297978
rect 316682 297922 316738 297978
rect 316806 297922 316862 297978
rect 316434 280294 316490 280350
rect 316558 280294 316614 280350
rect 316682 280294 316738 280350
rect 316806 280294 316862 280350
rect 316434 280170 316490 280226
rect 316558 280170 316614 280226
rect 316682 280170 316738 280226
rect 316806 280170 316862 280226
rect 316434 280046 316490 280102
rect 316558 280046 316614 280102
rect 316682 280046 316738 280102
rect 316806 280046 316862 280102
rect 316434 279922 316490 279978
rect 316558 279922 316614 279978
rect 316682 279922 316738 279978
rect 316806 279922 316862 279978
rect 316434 262294 316490 262350
rect 316558 262294 316614 262350
rect 316682 262294 316738 262350
rect 316806 262294 316862 262350
rect 316434 262170 316490 262226
rect 316558 262170 316614 262226
rect 316682 262170 316738 262226
rect 316806 262170 316862 262226
rect 316434 262046 316490 262102
rect 316558 262046 316614 262102
rect 316682 262046 316738 262102
rect 316806 262046 316862 262102
rect 316434 261922 316490 261978
rect 316558 261922 316614 261978
rect 316682 261922 316738 261978
rect 316806 261922 316862 261978
rect 316434 244294 316490 244350
rect 316558 244294 316614 244350
rect 316682 244294 316738 244350
rect 316806 244294 316862 244350
rect 316434 244170 316490 244226
rect 316558 244170 316614 244226
rect 316682 244170 316738 244226
rect 316806 244170 316862 244226
rect 316434 244046 316490 244102
rect 316558 244046 316614 244102
rect 316682 244046 316738 244102
rect 316806 244046 316862 244102
rect 316434 243922 316490 243978
rect 316558 243922 316614 243978
rect 316682 243922 316738 243978
rect 316806 243922 316862 243978
rect 316434 226294 316490 226350
rect 316558 226294 316614 226350
rect 316682 226294 316738 226350
rect 316806 226294 316862 226350
rect 316434 226170 316490 226226
rect 316558 226170 316614 226226
rect 316682 226170 316738 226226
rect 316806 226170 316862 226226
rect 316434 226046 316490 226102
rect 316558 226046 316614 226102
rect 316682 226046 316738 226102
rect 316806 226046 316862 226102
rect 316434 225922 316490 225978
rect 316558 225922 316614 225978
rect 316682 225922 316738 225978
rect 316806 225922 316862 225978
rect 316434 208294 316490 208350
rect 316558 208294 316614 208350
rect 316682 208294 316738 208350
rect 316806 208294 316862 208350
rect 316434 208170 316490 208226
rect 316558 208170 316614 208226
rect 316682 208170 316738 208226
rect 316806 208170 316862 208226
rect 316434 208046 316490 208102
rect 316558 208046 316614 208102
rect 316682 208046 316738 208102
rect 316806 208046 316862 208102
rect 316434 207922 316490 207978
rect 316558 207922 316614 207978
rect 316682 207922 316738 207978
rect 316806 207922 316862 207978
rect 316434 190294 316490 190350
rect 316558 190294 316614 190350
rect 316682 190294 316738 190350
rect 316806 190294 316862 190350
rect 316434 190170 316490 190226
rect 316558 190170 316614 190226
rect 316682 190170 316738 190226
rect 316806 190170 316862 190226
rect 316434 190046 316490 190102
rect 316558 190046 316614 190102
rect 316682 190046 316738 190102
rect 316806 190046 316862 190102
rect 316434 189922 316490 189978
rect 316558 189922 316614 189978
rect 316682 189922 316738 189978
rect 316806 189922 316862 189978
rect 316434 172294 316490 172350
rect 316558 172294 316614 172350
rect 316682 172294 316738 172350
rect 316806 172294 316862 172350
rect 316434 172170 316490 172226
rect 316558 172170 316614 172226
rect 316682 172170 316738 172226
rect 316806 172170 316862 172226
rect 316434 172046 316490 172102
rect 316558 172046 316614 172102
rect 316682 172046 316738 172102
rect 316806 172046 316862 172102
rect 316434 171922 316490 171978
rect 316558 171922 316614 171978
rect 316682 171922 316738 171978
rect 316806 171922 316862 171978
rect 343434 400294 343490 400350
rect 343558 400294 343614 400350
rect 343682 400294 343738 400350
rect 343806 400294 343862 400350
rect 343434 400170 343490 400226
rect 343558 400170 343614 400226
rect 343682 400170 343738 400226
rect 343806 400170 343862 400226
rect 343434 400046 343490 400102
rect 343558 400046 343614 400102
rect 343682 400046 343738 400102
rect 343806 400046 343862 400102
rect 343434 399922 343490 399978
rect 343558 399922 343614 399978
rect 343682 399922 343738 399978
rect 343806 399922 343862 399978
rect 343434 382294 343490 382350
rect 343558 382294 343614 382350
rect 343682 382294 343738 382350
rect 343806 382294 343862 382350
rect 343434 382170 343490 382226
rect 343558 382170 343614 382226
rect 343682 382170 343738 382226
rect 343806 382170 343862 382226
rect 343434 382046 343490 382102
rect 343558 382046 343614 382102
rect 343682 382046 343738 382102
rect 343806 382046 343862 382102
rect 343434 381922 343490 381978
rect 343558 381922 343614 381978
rect 343682 381922 343738 381978
rect 343806 381922 343862 381978
rect 343434 364294 343490 364350
rect 343558 364294 343614 364350
rect 343682 364294 343738 364350
rect 343806 364294 343862 364350
rect 343434 364170 343490 364226
rect 343558 364170 343614 364226
rect 343682 364170 343738 364226
rect 343806 364170 343862 364226
rect 343434 364046 343490 364102
rect 343558 364046 343614 364102
rect 343682 364046 343738 364102
rect 343806 364046 343862 364102
rect 343434 363922 343490 363978
rect 343558 363922 343614 363978
rect 343682 363922 343738 363978
rect 343806 363922 343862 363978
rect 343434 346294 343490 346350
rect 343558 346294 343614 346350
rect 343682 346294 343738 346350
rect 343806 346294 343862 346350
rect 343434 346170 343490 346226
rect 343558 346170 343614 346226
rect 343682 346170 343738 346226
rect 343806 346170 343862 346226
rect 343434 346046 343490 346102
rect 343558 346046 343614 346102
rect 343682 346046 343738 346102
rect 343806 346046 343862 346102
rect 343434 345922 343490 345978
rect 343558 345922 343614 345978
rect 343682 345922 343738 345978
rect 343806 345922 343862 345978
rect 343434 328294 343490 328350
rect 343558 328294 343614 328350
rect 343682 328294 343738 328350
rect 343806 328294 343862 328350
rect 343434 328170 343490 328226
rect 343558 328170 343614 328226
rect 343682 328170 343738 328226
rect 343806 328170 343862 328226
rect 343434 328046 343490 328102
rect 343558 328046 343614 328102
rect 343682 328046 343738 328102
rect 343806 328046 343862 328102
rect 343434 327922 343490 327978
rect 343558 327922 343614 327978
rect 343682 327922 343738 327978
rect 343806 327922 343862 327978
rect 343434 310294 343490 310350
rect 343558 310294 343614 310350
rect 343682 310294 343738 310350
rect 343806 310294 343862 310350
rect 343434 310170 343490 310226
rect 343558 310170 343614 310226
rect 343682 310170 343738 310226
rect 343806 310170 343862 310226
rect 343434 310046 343490 310102
rect 343558 310046 343614 310102
rect 343682 310046 343738 310102
rect 343806 310046 343862 310102
rect 343434 309922 343490 309978
rect 343558 309922 343614 309978
rect 343682 309922 343738 309978
rect 343806 309922 343862 309978
rect 343434 292294 343490 292350
rect 343558 292294 343614 292350
rect 343682 292294 343738 292350
rect 343806 292294 343862 292350
rect 343434 292170 343490 292226
rect 343558 292170 343614 292226
rect 343682 292170 343738 292226
rect 343806 292170 343862 292226
rect 343434 292046 343490 292102
rect 343558 292046 343614 292102
rect 343682 292046 343738 292102
rect 343806 292046 343862 292102
rect 343434 291922 343490 291978
rect 343558 291922 343614 291978
rect 343682 291922 343738 291978
rect 343806 291922 343862 291978
rect 343434 274294 343490 274350
rect 343558 274294 343614 274350
rect 343682 274294 343738 274350
rect 343806 274294 343862 274350
rect 343434 274170 343490 274226
rect 343558 274170 343614 274226
rect 343682 274170 343738 274226
rect 343806 274170 343862 274226
rect 343434 274046 343490 274102
rect 343558 274046 343614 274102
rect 343682 274046 343738 274102
rect 343806 274046 343862 274102
rect 343434 273922 343490 273978
rect 343558 273922 343614 273978
rect 343682 273922 343738 273978
rect 343806 273922 343862 273978
rect 343434 256294 343490 256350
rect 343558 256294 343614 256350
rect 343682 256294 343738 256350
rect 343806 256294 343862 256350
rect 343434 256170 343490 256226
rect 343558 256170 343614 256226
rect 343682 256170 343738 256226
rect 343806 256170 343862 256226
rect 343434 256046 343490 256102
rect 343558 256046 343614 256102
rect 343682 256046 343738 256102
rect 343806 256046 343862 256102
rect 343434 255922 343490 255978
rect 343558 255922 343614 255978
rect 343682 255922 343738 255978
rect 343806 255922 343862 255978
rect 343434 238294 343490 238350
rect 343558 238294 343614 238350
rect 343682 238294 343738 238350
rect 343806 238294 343862 238350
rect 343434 238170 343490 238226
rect 343558 238170 343614 238226
rect 343682 238170 343738 238226
rect 343806 238170 343862 238226
rect 343434 238046 343490 238102
rect 343558 238046 343614 238102
rect 343682 238046 343738 238102
rect 343806 238046 343862 238102
rect 343434 237922 343490 237978
rect 343558 237922 343614 237978
rect 343682 237922 343738 237978
rect 343806 237922 343862 237978
rect 343434 220294 343490 220350
rect 343558 220294 343614 220350
rect 343682 220294 343738 220350
rect 343806 220294 343862 220350
rect 343434 220170 343490 220226
rect 343558 220170 343614 220226
rect 343682 220170 343738 220226
rect 343806 220170 343862 220226
rect 343434 220046 343490 220102
rect 343558 220046 343614 220102
rect 343682 220046 343738 220102
rect 343806 220046 343862 220102
rect 343434 219922 343490 219978
rect 343558 219922 343614 219978
rect 343682 219922 343738 219978
rect 343806 219922 343862 219978
rect 343434 202294 343490 202350
rect 343558 202294 343614 202350
rect 343682 202294 343738 202350
rect 343806 202294 343862 202350
rect 343434 202170 343490 202226
rect 343558 202170 343614 202226
rect 343682 202170 343738 202226
rect 343806 202170 343862 202226
rect 343434 202046 343490 202102
rect 343558 202046 343614 202102
rect 343682 202046 343738 202102
rect 343806 202046 343862 202102
rect 343434 201922 343490 201978
rect 343558 201922 343614 201978
rect 343682 201922 343738 201978
rect 343806 201922 343862 201978
rect 343434 184294 343490 184350
rect 343558 184294 343614 184350
rect 343682 184294 343738 184350
rect 343806 184294 343862 184350
rect 343434 184170 343490 184226
rect 343558 184170 343614 184226
rect 343682 184170 343738 184226
rect 343806 184170 343862 184226
rect 343434 184046 343490 184102
rect 343558 184046 343614 184102
rect 343682 184046 343738 184102
rect 343806 184046 343862 184102
rect 343434 183922 343490 183978
rect 343558 183922 343614 183978
rect 343682 183922 343738 183978
rect 343806 183922 343862 183978
rect 343434 166294 343490 166350
rect 343558 166294 343614 166350
rect 343682 166294 343738 166350
rect 343806 166294 343862 166350
rect 343434 166170 343490 166226
rect 343558 166170 343614 166226
rect 343682 166170 343738 166226
rect 343806 166170 343862 166226
rect 343434 166046 343490 166102
rect 343558 166046 343614 166102
rect 343682 166046 343738 166102
rect 343806 166046 343862 166102
rect 343434 165922 343490 165978
rect 343558 165922 343614 165978
rect 343682 165922 343738 165978
rect 343806 165922 343862 165978
rect 316434 154294 316490 154350
rect 316558 154294 316614 154350
rect 316682 154294 316738 154350
rect 316806 154294 316862 154350
rect 316434 154170 316490 154226
rect 316558 154170 316614 154226
rect 316682 154170 316738 154226
rect 316806 154170 316862 154226
rect 316434 154046 316490 154102
rect 316558 154046 316614 154102
rect 316682 154046 316738 154102
rect 316806 154046 316862 154102
rect 316434 153922 316490 153978
rect 316558 153922 316614 153978
rect 316682 153922 316738 153978
rect 316806 153922 316862 153978
rect 314636 141002 314692 141058
rect 312714 130294 312770 130350
rect 312838 130294 312894 130350
rect 312962 130294 313018 130350
rect 313086 130294 313142 130350
rect 312714 130170 312770 130226
rect 312838 130170 312894 130226
rect 312962 130170 313018 130226
rect 313086 130170 313142 130226
rect 312714 130046 312770 130102
rect 312838 130046 312894 130102
rect 312962 130046 313018 130102
rect 313086 130046 313142 130102
rect 312714 129922 312770 129978
rect 312838 129922 312894 129978
rect 312962 129922 313018 129978
rect 313086 129922 313142 129978
rect 312714 112294 312770 112350
rect 312838 112294 312894 112350
rect 312962 112294 313018 112350
rect 313086 112294 313142 112350
rect 312714 112170 312770 112226
rect 312838 112170 312894 112226
rect 312962 112170 313018 112226
rect 313086 112170 313142 112226
rect 312714 112046 312770 112102
rect 312838 112046 312894 112102
rect 312962 112046 313018 112102
rect 313086 112046 313142 112102
rect 312714 111922 312770 111978
rect 312838 111922 312894 111978
rect 312962 111922 313018 111978
rect 313086 111922 313142 111978
rect 312714 94294 312770 94350
rect 312838 94294 312894 94350
rect 312962 94294 313018 94350
rect 313086 94294 313142 94350
rect 312714 94170 312770 94226
rect 312838 94170 312894 94226
rect 312962 94170 313018 94226
rect 313086 94170 313142 94226
rect 312714 94046 312770 94102
rect 312838 94046 312894 94102
rect 312962 94046 313018 94102
rect 313086 94046 313142 94102
rect 312714 93922 312770 93978
rect 312838 93922 312894 93978
rect 312962 93922 313018 93978
rect 313086 93922 313142 93978
rect 312714 76294 312770 76350
rect 312838 76294 312894 76350
rect 312962 76294 313018 76350
rect 313086 76294 313142 76350
rect 312714 76170 312770 76226
rect 312838 76170 312894 76226
rect 312962 76170 313018 76226
rect 313086 76170 313142 76226
rect 312714 76046 312770 76102
rect 312838 76046 312894 76102
rect 312962 76046 313018 76102
rect 313086 76046 313142 76102
rect 312714 75922 312770 75978
rect 312838 75922 312894 75978
rect 312962 75922 313018 75978
rect 313086 75922 313142 75978
rect 312714 58294 312770 58350
rect 312838 58294 312894 58350
rect 312962 58294 313018 58350
rect 313086 58294 313142 58350
rect 312714 58170 312770 58226
rect 312838 58170 312894 58226
rect 312962 58170 313018 58226
rect 313086 58170 313142 58226
rect 312714 58046 312770 58102
rect 312838 58046 312894 58102
rect 312962 58046 313018 58102
rect 313086 58046 313142 58102
rect 312714 57922 312770 57978
rect 312838 57922 312894 57978
rect 312962 57922 313018 57978
rect 313086 57922 313142 57978
rect 312714 40294 312770 40350
rect 312838 40294 312894 40350
rect 312962 40294 313018 40350
rect 313086 40294 313142 40350
rect 312714 40170 312770 40226
rect 312838 40170 312894 40226
rect 312962 40170 313018 40226
rect 313086 40170 313142 40226
rect 312714 40046 312770 40102
rect 312838 40046 312894 40102
rect 312962 40046 313018 40102
rect 313086 40046 313142 40102
rect 312714 39922 312770 39978
rect 312838 39922 312894 39978
rect 312962 39922 313018 39978
rect 313086 39922 313142 39978
rect 312714 22294 312770 22350
rect 312838 22294 312894 22350
rect 312962 22294 313018 22350
rect 313086 22294 313142 22350
rect 312714 22170 312770 22226
rect 312838 22170 312894 22226
rect 312962 22170 313018 22226
rect 313086 22170 313142 22226
rect 312714 22046 312770 22102
rect 312838 22046 312894 22102
rect 312962 22046 313018 22102
rect 313086 22046 313142 22102
rect 312714 21922 312770 21978
rect 312838 21922 312894 21978
rect 312962 21922 313018 21978
rect 313086 21922 313142 21978
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 285714 -1176 285770 -1120
rect 285838 -1176 285894 -1120
rect 285962 -1176 286018 -1120
rect 286086 -1176 286142 -1120
rect 285714 -1300 285770 -1244
rect 285838 -1300 285894 -1244
rect 285962 -1300 286018 -1244
rect 286086 -1300 286142 -1244
rect 285714 -1424 285770 -1368
rect 285838 -1424 285894 -1368
rect 285962 -1424 286018 -1368
rect 286086 -1424 286142 -1368
rect 285714 -1548 285770 -1492
rect 285838 -1548 285894 -1492
rect 285962 -1548 286018 -1492
rect 286086 -1548 286142 -1492
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 319228 141902 319284 141958
rect 316434 136294 316490 136350
rect 316558 136294 316614 136350
rect 316682 136294 316738 136350
rect 316806 136294 316862 136350
rect 316434 136170 316490 136226
rect 316558 136170 316614 136226
rect 316682 136170 316738 136226
rect 316806 136170 316862 136226
rect 316434 136046 316490 136102
rect 316558 136046 316614 136102
rect 316682 136046 316738 136102
rect 316806 136046 316862 136102
rect 316434 135922 316490 135978
rect 316558 135922 316614 135978
rect 316682 135922 316738 135978
rect 316806 135922 316862 135978
rect 316434 118294 316490 118350
rect 316558 118294 316614 118350
rect 316682 118294 316738 118350
rect 316806 118294 316862 118350
rect 316434 118170 316490 118226
rect 316558 118170 316614 118226
rect 316682 118170 316738 118226
rect 316806 118170 316862 118226
rect 316434 118046 316490 118102
rect 316558 118046 316614 118102
rect 316682 118046 316738 118102
rect 316806 118046 316862 118102
rect 316434 117922 316490 117978
rect 316558 117922 316614 117978
rect 316682 117922 316738 117978
rect 316806 117922 316862 117978
rect 316434 100294 316490 100350
rect 316558 100294 316614 100350
rect 316682 100294 316738 100350
rect 316806 100294 316862 100350
rect 316434 100170 316490 100226
rect 316558 100170 316614 100226
rect 316682 100170 316738 100226
rect 316806 100170 316862 100226
rect 316434 100046 316490 100102
rect 316558 100046 316614 100102
rect 316682 100046 316738 100102
rect 316806 100046 316862 100102
rect 316434 99922 316490 99978
rect 316558 99922 316614 99978
rect 316682 99922 316738 99978
rect 316806 99922 316862 99978
rect 316434 82294 316490 82350
rect 316558 82294 316614 82350
rect 316682 82294 316738 82350
rect 316806 82294 316862 82350
rect 316434 82170 316490 82226
rect 316558 82170 316614 82226
rect 316682 82170 316738 82226
rect 316806 82170 316862 82226
rect 316434 82046 316490 82102
rect 316558 82046 316614 82102
rect 316682 82046 316738 82102
rect 316806 82046 316862 82102
rect 316434 81922 316490 81978
rect 316558 81922 316614 81978
rect 316682 81922 316738 81978
rect 316806 81922 316862 81978
rect 316434 64294 316490 64350
rect 316558 64294 316614 64350
rect 316682 64294 316738 64350
rect 316806 64294 316862 64350
rect 316434 64170 316490 64226
rect 316558 64170 316614 64226
rect 316682 64170 316738 64226
rect 316806 64170 316862 64226
rect 316434 64046 316490 64102
rect 316558 64046 316614 64102
rect 316682 64046 316738 64102
rect 316806 64046 316862 64102
rect 316434 63922 316490 63978
rect 316558 63922 316614 63978
rect 316682 63922 316738 63978
rect 316806 63922 316862 63978
rect 316434 46294 316490 46350
rect 316558 46294 316614 46350
rect 316682 46294 316738 46350
rect 316806 46294 316862 46350
rect 316434 46170 316490 46226
rect 316558 46170 316614 46226
rect 316682 46170 316738 46226
rect 316806 46170 316862 46226
rect 316434 46046 316490 46102
rect 316558 46046 316614 46102
rect 316682 46046 316738 46102
rect 316806 46046 316862 46102
rect 316434 45922 316490 45978
rect 316558 45922 316614 45978
rect 316682 45922 316738 45978
rect 316806 45922 316862 45978
rect 316434 28294 316490 28350
rect 316558 28294 316614 28350
rect 316682 28294 316738 28350
rect 316806 28294 316862 28350
rect 316434 28170 316490 28226
rect 316558 28170 316614 28226
rect 316682 28170 316738 28226
rect 316806 28170 316862 28226
rect 316434 28046 316490 28102
rect 316558 28046 316614 28102
rect 316682 28046 316738 28102
rect 316806 28046 316862 28102
rect 316434 27922 316490 27978
rect 316558 27922 316614 27978
rect 316682 27922 316738 27978
rect 316806 27922 316862 27978
rect 316434 10294 316490 10350
rect 316558 10294 316614 10350
rect 316682 10294 316738 10350
rect 316806 10294 316862 10350
rect 316434 10170 316490 10226
rect 316558 10170 316614 10226
rect 316682 10170 316738 10226
rect 316806 10170 316862 10226
rect 316434 10046 316490 10102
rect 316558 10046 316614 10102
rect 316682 10046 316738 10102
rect 316806 10046 316862 10102
rect 316434 9922 316490 9978
rect 316558 9922 316614 9978
rect 316682 9922 316738 9978
rect 316806 9922 316862 9978
rect 343434 148294 343490 148350
rect 343558 148294 343614 148350
rect 343682 148294 343738 148350
rect 343806 148294 343862 148350
rect 343434 148170 343490 148226
rect 343558 148170 343614 148226
rect 343682 148170 343738 148226
rect 343806 148170 343862 148226
rect 343434 148046 343490 148102
rect 343558 148046 343614 148102
rect 343682 148046 343738 148102
rect 343806 148046 343862 148102
rect 343434 147922 343490 147978
rect 343558 147922 343614 147978
rect 343682 147922 343738 147978
rect 343806 147922 343862 147978
rect 330876 141902 330932 141958
rect 333452 141002 333508 141058
rect 340956 140822 341012 140878
rect 347154 388294 347210 388350
rect 347278 388294 347334 388350
rect 347402 388294 347458 388350
rect 347526 388294 347582 388350
rect 347154 388170 347210 388226
rect 347278 388170 347334 388226
rect 347402 388170 347458 388226
rect 347526 388170 347582 388226
rect 347154 388046 347210 388102
rect 347278 388046 347334 388102
rect 347402 388046 347458 388102
rect 347526 388046 347582 388102
rect 347154 387922 347210 387978
rect 347278 387922 347334 387978
rect 347402 387922 347458 387978
rect 347526 387922 347582 387978
rect 347154 370294 347210 370350
rect 347278 370294 347334 370350
rect 347402 370294 347458 370350
rect 347526 370294 347582 370350
rect 347154 370170 347210 370226
rect 347278 370170 347334 370226
rect 347402 370170 347458 370226
rect 347526 370170 347582 370226
rect 347154 370046 347210 370102
rect 347278 370046 347334 370102
rect 347402 370046 347458 370102
rect 347526 370046 347582 370102
rect 347154 369922 347210 369978
rect 347278 369922 347334 369978
rect 347402 369922 347458 369978
rect 347526 369922 347582 369978
rect 347154 352294 347210 352350
rect 347278 352294 347334 352350
rect 347402 352294 347458 352350
rect 347526 352294 347582 352350
rect 347154 352170 347210 352226
rect 347278 352170 347334 352226
rect 347402 352170 347458 352226
rect 347526 352170 347582 352226
rect 347154 352046 347210 352102
rect 347278 352046 347334 352102
rect 347402 352046 347458 352102
rect 347526 352046 347582 352102
rect 347154 351922 347210 351978
rect 347278 351922 347334 351978
rect 347402 351922 347458 351978
rect 347526 351922 347582 351978
rect 374154 400294 374210 400350
rect 374278 400294 374334 400350
rect 374402 400294 374458 400350
rect 374526 400294 374582 400350
rect 374154 400170 374210 400226
rect 374278 400170 374334 400226
rect 374402 400170 374458 400226
rect 374526 400170 374582 400226
rect 374154 400046 374210 400102
rect 374278 400046 374334 400102
rect 374402 400046 374458 400102
rect 374526 400046 374582 400102
rect 374154 399922 374210 399978
rect 374278 399922 374334 399978
rect 374402 399922 374458 399978
rect 374526 399922 374582 399978
rect 374154 382294 374210 382350
rect 374278 382294 374334 382350
rect 374402 382294 374458 382350
rect 374526 382294 374582 382350
rect 374154 382170 374210 382226
rect 374278 382170 374334 382226
rect 374402 382170 374458 382226
rect 374526 382170 374582 382226
rect 374154 382046 374210 382102
rect 374278 382046 374334 382102
rect 374402 382046 374458 382102
rect 374526 382046 374582 382102
rect 374154 381922 374210 381978
rect 374278 381922 374334 381978
rect 374402 381922 374458 381978
rect 374526 381922 374582 381978
rect 374154 364294 374210 364350
rect 374278 364294 374334 364350
rect 374402 364294 374458 364350
rect 374526 364294 374582 364350
rect 374154 364170 374210 364226
rect 374278 364170 374334 364226
rect 374402 364170 374458 364226
rect 374526 364170 374582 364226
rect 374154 364046 374210 364102
rect 374278 364046 374334 364102
rect 374402 364046 374458 364102
rect 374526 364046 374582 364102
rect 374154 363922 374210 363978
rect 374278 363922 374334 363978
rect 374402 363922 374458 363978
rect 374526 363922 374582 363978
rect 347154 334294 347210 334350
rect 347278 334294 347334 334350
rect 347402 334294 347458 334350
rect 347526 334294 347582 334350
rect 347154 334170 347210 334226
rect 347278 334170 347334 334226
rect 347402 334170 347458 334226
rect 347526 334170 347582 334226
rect 347154 334046 347210 334102
rect 347278 334046 347334 334102
rect 347402 334046 347458 334102
rect 347526 334046 347582 334102
rect 347154 333922 347210 333978
rect 347278 333922 347334 333978
rect 347402 333922 347458 333978
rect 347526 333922 347582 333978
rect 355292 349442 355348 349498
rect 351932 330002 351988 330058
rect 347154 316294 347210 316350
rect 347278 316294 347334 316350
rect 347402 316294 347458 316350
rect 347526 316294 347582 316350
rect 347154 316170 347210 316226
rect 347278 316170 347334 316226
rect 347402 316170 347458 316226
rect 347526 316170 347582 316226
rect 347154 316046 347210 316102
rect 347278 316046 347334 316102
rect 347402 316046 347458 316102
rect 347526 316046 347582 316102
rect 347154 315922 347210 315978
rect 347278 315922 347334 315978
rect 347402 315922 347458 315978
rect 347526 315922 347582 315978
rect 347154 298294 347210 298350
rect 347278 298294 347334 298350
rect 347402 298294 347458 298350
rect 347526 298294 347582 298350
rect 347154 298170 347210 298226
rect 347278 298170 347334 298226
rect 347402 298170 347458 298226
rect 347526 298170 347582 298226
rect 347154 298046 347210 298102
rect 347278 298046 347334 298102
rect 347402 298046 347458 298102
rect 347526 298046 347582 298102
rect 347154 297922 347210 297978
rect 347278 297922 347334 297978
rect 347402 297922 347458 297978
rect 347526 297922 347582 297978
rect 347154 280294 347210 280350
rect 347278 280294 347334 280350
rect 347402 280294 347458 280350
rect 347526 280294 347582 280350
rect 347154 280170 347210 280226
rect 347278 280170 347334 280226
rect 347402 280170 347458 280226
rect 347526 280170 347582 280226
rect 347154 280046 347210 280102
rect 347278 280046 347334 280102
rect 347402 280046 347458 280102
rect 347526 280046 347582 280102
rect 347154 279922 347210 279978
rect 347278 279922 347334 279978
rect 347402 279922 347458 279978
rect 347526 279922 347582 279978
rect 347154 262294 347210 262350
rect 347278 262294 347334 262350
rect 347402 262294 347458 262350
rect 347526 262294 347582 262350
rect 347154 262170 347210 262226
rect 347278 262170 347334 262226
rect 347402 262170 347458 262226
rect 347526 262170 347582 262226
rect 347154 262046 347210 262102
rect 347278 262046 347334 262102
rect 347402 262046 347458 262102
rect 347526 262046 347582 262102
rect 347154 261922 347210 261978
rect 347278 261922 347334 261978
rect 347402 261922 347458 261978
rect 347526 261922 347582 261978
rect 347154 244294 347210 244350
rect 347278 244294 347334 244350
rect 347402 244294 347458 244350
rect 347526 244294 347582 244350
rect 347154 244170 347210 244226
rect 347278 244170 347334 244226
rect 347402 244170 347458 244226
rect 347526 244170 347582 244226
rect 347154 244046 347210 244102
rect 347278 244046 347334 244102
rect 347402 244046 347458 244102
rect 347526 244046 347582 244102
rect 347154 243922 347210 243978
rect 347278 243922 347334 243978
rect 347402 243922 347458 243978
rect 347526 243922 347582 243978
rect 347154 226294 347210 226350
rect 347278 226294 347334 226350
rect 347402 226294 347458 226350
rect 347526 226294 347582 226350
rect 347154 226170 347210 226226
rect 347278 226170 347334 226226
rect 347402 226170 347458 226226
rect 347526 226170 347582 226226
rect 347154 226046 347210 226102
rect 347278 226046 347334 226102
rect 347402 226046 347458 226102
rect 347526 226046 347582 226102
rect 347154 225922 347210 225978
rect 347278 225922 347334 225978
rect 347402 225922 347458 225978
rect 347526 225922 347582 225978
rect 347154 208294 347210 208350
rect 347278 208294 347334 208350
rect 347402 208294 347458 208350
rect 347526 208294 347582 208350
rect 347154 208170 347210 208226
rect 347278 208170 347334 208226
rect 347402 208170 347458 208226
rect 347526 208170 347582 208226
rect 347154 208046 347210 208102
rect 347278 208046 347334 208102
rect 347402 208046 347458 208102
rect 347526 208046 347582 208102
rect 347154 207922 347210 207978
rect 347278 207922 347334 207978
rect 347402 207922 347458 207978
rect 347526 207922 347582 207978
rect 347154 190294 347210 190350
rect 347278 190294 347334 190350
rect 347402 190294 347458 190350
rect 347526 190294 347582 190350
rect 347154 190170 347210 190226
rect 347278 190170 347334 190226
rect 347402 190170 347458 190226
rect 347526 190170 347582 190226
rect 347154 190046 347210 190102
rect 347278 190046 347334 190102
rect 347402 190046 347458 190102
rect 347526 190046 347582 190102
rect 347154 189922 347210 189978
rect 347278 189922 347334 189978
rect 347402 189922 347458 189978
rect 347526 189922 347582 189978
rect 347154 172294 347210 172350
rect 347278 172294 347334 172350
rect 347402 172294 347458 172350
rect 347526 172294 347582 172350
rect 347154 172170 347210 172226
rect 347278 172170 347334 172226
rect 347402 172170 347458 172226
rect 347526 172170 347582 172226
rect 347154 172046 347210 172102
rect 347278 172046 347334 172102
rect 347402 172046 347458 172102
rect 347526 172046 347582 172102
rect 347154 171922 347210 171978
rect 347278 171922 347334 171978
rect 347402 171922 347458 171978
rect 347526 171922 347582 171978
rect 347154 154294 347210 154350
rect 347278 154294 347334 154350
rect 347402 154294 347458 154350
rect 347526 154294 347582 154350
rect 347154 154170 347210 154226
rect 347278 154170 347334 154226
rect 347402 154170 347458 154226
rect 347526 154170 347582 154226
rect 347154 154046 347210 154102
rect 347278 154046 347334 154102
rect 347402 154046 347458 154102
rect 347526 154046 347582 154102
rect 347154 153922 347210 153978
rect 347278 153922 347334 153978
rect 347402 153922 347458 153978
rect 347526 153922 347582 153978
rect 344652 142100 344708 142138
rect 344652 142082 344708 142100
rect 348572 319922 348628 319978
rect 343434 130294 343490 130350
rect 343558 130294 343614 130350
rect 343682 130294 343738 130350
rect 343806 130294 343862 130350
rect 343434 130170 343490 130226
rect 343558 130170 343614 130226
rect 343682 130170 343738 130226
rect 343806 130170 343862 130226
rect 343434 130046 343490 130102
rect 343558 130046 343614 130102
rect 343682 130046 343738 130102
rect 343806 130046 343862 130102
rect 343434 129922 343490 129978
rect 343558 129922 343614 129978
rect 343682 129922 343738 129978
rect 343806 129922 343862 129978
rect 345812 130294 345868 130350
rect 345936 130294 345992 130350
rect 346060 130294 346116 130350
rect 346184 130294 346240 130350
rect 345812 130170 345868 130226
rect 345936 130170 345992 130226
rect 346060 130170 346116 130226
rect 346184 130170 346240 130226
rect 345812 130046 345868 130102
rect 345936 130046 345992 130102
rect 346060 130046 346116 130102
rect 346184 130046 346240 130102
rect 345812 129922 345868 129978
rect 345936 129922 345992 129978
rect 346060 129922 346116 129978
rect 346184 129922 346240 129978
rect 346612 118294 346668 118350
rect 346736 118294 346792 118350
rect 346860 118294 346916 118350
rect 346984 118294 347040 118350
rect 346612 118170 346668 118226
rect 346736 118170 346792 118226
rect 346860 118170 346916 118226
rect 346984 118170 347040 118226
rect 346612 118046 346668 118102
rect 346736 118046 346792 118102
rect 346860 118046 346916 118102
rect 346984 118046 347040 118102
rect 346612 117922 346668 117978
rect 346736 117922 346792 117978
rect 346860 117922 346916 117978
rect 346984 117922 347040 117978
rect 343434 112294 343490 112350
rect 343558 112294 343614 112350
rect 343682 112294 343738 112350
rect 343806 112294 343862 112350
rect 343434 112170 343490 112226
rect 343558 112170 343614 112226
rect 343682 112170 343738 112226
rect 343806 112170 343862 112226
rect 343434 112046 343490 112102
rect 343558 112046 343614 112102
rect 343682 112046 343738 112102
rect 343806 112046 343862 112102
rect 343434 111922 343490 111978
rect 343558 111922 343614 111978
rect 343682 111922 343738 111978
rect 343806 111922 343862 111978
rect 345812 112294 345868 112350
rect 345936 112294 345992 112350
rect 346060 112294 346116 112350
rect 346184 112294 346240 112350
rect 345812 112170 345868 112226
rect 345936 112170 345992 112226
rect 346060 112170 346116 112226
rect 346184 112170 346240 112226
rect 345812 112046 345868 112102
rect 345936 112046 345992 112102
rect 346060 112046 346116 112102
rect 346184 112046 346240 112102
rect 345812 111922 345868 111978
rect 345936 111922 345992 111978
rect 346060 111922 346116 111978
rect 346184 111922 346240 111978
rect 346612 100294 346668 100350
rect 346736 100294 346792 100350
rect 346860 100294 346916 100350
rect 346984 100294 347040 100350
rect 346612 100170 346668 100226
rect 346736 100170 346792 100226
rect 346860 100170 346916 100226
rect 346984 100170 347040 100226
rect 346612 100046 346668 100102
rect 346736 100046 346792 100102
rect 346860 100046 346916 100102
rect 346984 100046 347040 100102
rect 346612 99922 346668 99978
rect 346736 99922 346792 99978
rect 346860 99922 346916 99978
rect 346984 99922 347040 99978
rect 343434 94294 343490 94350
rect 343558 94294 343614 94350
rect 343682 94294 343738 94350
rect 343806 94294 343862 94350
rect 343434 94170 343490 94226
rect 343558 94170 343614 94226
rect 343682 94170 343738 94226
rect 343806 94170 343862 94226
rect 343434 94046 343490 94102
rect 343558 94046 343614 94102
rect 343682 94046 343738 94102
rect 343806 94046 343862 94102
rect 343434 93922 343490 93978
rect 343558 93922 343614 93978
rect 343682 93922 343738 93978
rect 343806 93922 343862 93978
rect 345812 94294 345868 94350
rect 345936 94294 345992 94350
rect 346060 94294 346116 94350
rect 346184 94294 346240 94350
rect 345812 94170 345868 94226
rect 345936 94170 345992 94226
rect 346060 94170 346116 94226
rect 346184 94170 346240 94226
rect 345812 94046 345868 94102
rect 345936 94046 345992 94102
rect 346060 94046 346116 94102
rect 346184 94046 346240 94102
rect 345812 93922 345868 93978
rect 345936 93922 345992 93978
rect 346060 93922 346116 93978
rect 346184 93922 346240 93978
rect 346612 82294 346668 82350
rect 346736 82294 346792 82350
rect 346860 82294 346916 82350
rect 346984 82294 347040 82350
rect 346612 82170 346668 82226
rect 346736 82170 346792 82226
rect 346860 82170 346916 82226
rect 346984 82170 347040 82226
rect 346612 82046 346668 82102
rect 346736 82046 346792 82102
rect 346860 82046 346916 82102
rect 346984 82046 347040 82102
rect 346612 81922 346668 81978
rect 346736 81922 346792 81978
rect 346860 81922 346916 81978
rect 346984 81922 347040 81978
rect 343434 76294 343490 76350
rect 343558 76294 343614 76350
rect 343682 76294 343738 76350
rect 343806 76294 343862 76350
rect 343434 76170 343490 76226
rect 343558 76170 343614 76226
rect 343682 76170 343738 76226
rect 343806 76170 343862 76226
rect 343434 76046 343490 76102
rect 343558 76046 343614 76102
rect 343682 76046 343738 76102
rect 343806 76046 343862 76102
rect 343434 75922 343490 75978
rect 343558 75922 343614 75978
rect 343682 75922 343738 75978
rect 343806 75922 343862 75978
rect 345812 76294 345868 76350
rect 345936 76294 345992 76350
rect 346060 76294 346116 76350
rect 346184 76294 346240 76350
rect 345812 76170 345868 76226
rect 345936 76170 345992 76226
rect 346060 76170 346116 76226
rect 346184 76170 346240 76226
rect 345812 76046 345868 76102
rect 345936 76046 345992 76102
rect 346060 76046 346116 76102
rect 346184 76046 346240 76102
rect 345812 75922 345868 75978
rect 345936 75922 345992 75978
rect 346060 75922 346116 75978
rect 346184 75922 346240 75978
rect 346612 64294 346668 64350
rect 346736 64294 346792 64350
rect 346860 64294 346916 64350
rect 346984 64294 347040 64350
rect 346612 64170 346668 64226
rect 346736 64170 346792 64226
rect 346860 64170 346916 64226
rect 346984 64170 347040 64226
rect 346612 64046 346668 64102
rect 346736 64046 346792 64102
rect 346860 64046 346916 64102
rect 346984 64046 347040 64102
rect 346612 63922 346668 63978
rect 346736 63922 346792 63978
rect 346860 63922 346916 63978
rect 346984 63922 347040 63978
rect 343434 58294 343490 58350
rect 343558 58294 343614 58350
rect 343682 58294 343738 58350
rect 343806 58294 343862 58350
rect 343434 58170 343490 58226
rect 343558 58170 343614 58226
rect 343682 58170 343738 58226
rect 343806 58170 343862 58226
rect 343434 58046 343490 58102
rect 343558 58046 343614 58102
rect 343682 58046 343738 58102
rect 343806 58046 343862 58102
rect 343434 57922 343490 57978
rect 343558 57922 343614 57978
rect 343682 57922 343738 57978
rect 343806 57922 343862 57978
rect 345812 58294 345868 58350
rect 345936 58294 345992 58350
rect 346060 58294 346116 58350
rect 346184 58294 346240 58350
rect 345812 58170 345868 58226
rect 345936 58170 345992 58226
rect 346060 58170 346116 58226
rect 346184 58170 346240 58226
rect 345812 58046 345868 58102
rect 345936 58046 345992 58102
rect 346060 58046 346116 58102
rect 346184 58046 346240 58102
rect 345812 57922 345868 57978
rect 345936 57922 345992 57978
rect 346060 57922 346116 57978
rect 346184 57922 346240 57978
rect 346612 46294 346668 46350
rect 346736 46294 346792 46350
rect 346860 46294 346916 46350
rect 346984 46294 347040 46350
rect 346612 46170 346668 46226
rect 346736 46170 346792 46226
rect 346860 46170 346916 46226
rect 346984 46170 347040 46226
rect 346612 46046 346668 46102
rect 346736 46046 346792 46102
rect 346860 46046 346916 46102
rect 346984 46046 347040 46102
rect 346612 45922 346668 45978
rect 346736 45922 346792 45978
rect 346860 45922 346916 45978
rect 346984 45922 347040 45978
rect 343434 40294 343490 40350
rect 343558 40294 343614 40350
rect 343682 40294 343738 40350
rect 343806 40294 343862 40350
rect 343434 40170 343490 40226
rect 343558 40170 343614 40226
rect 343682 40170 343738 40226
rect 343806 40170 343862 40226
rect 343434 40046 343490 40102
rect 343558 40046 343614 40102
rect 343682 40046 343738 40102
rect 343806 40046 343862 40102
rect 343434 39922 343490 39978
rect 343558 39922 343614 39978
rect 343682 39922 343738 39978
rect 343806 39922 343862 39978
rect 343434 22294 343490 22350
rect 343558 22294 343614 22350
rect 343682 22294 343738 22350
rect 343806 22294 343862 22350
rect 343434 22170 343490 22226
rect 343558 22170 343614 22226
rect 343682 22170 343738 22226
rect 343806 22170 343862 22226
rect 343434 22046 343490 22102
rect 343558 22046 343614 22102
rect 343682 22046 343738 22102
rect 343806 22046 343862 22102
rect 343434 21922 343490 21978
rect 343558 21922 343614 21978
rect 343682 21922 343738 21978
rect 343806 21922 343862 21978
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 316434 -1176 316490 -1120
rect 316558 -1176 316614 -1120
rect 316682 -1176 316738 -1120
rect 316806 -1176 316862 -1120
rect 316434 -1300 316490 -1244
rect 316558 -1300 316614 -1244
rect 316682 -1300 316738 -1244
rect 316806 -1300 316862 -1244
rect 316434 -1424 316490 -1368
rect 316558 -1424 316614 -1368
rect 316682 -1424 316738 -1368
rect 316806 -1424 316862 -1368
rect 316434 -1548 316490 -1492
rect 316558 -1548 316614 -1492
rect 316682 -1548 316738 -1492
rect 316806 -1548 316862 -1492
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 347154 28294 347210 28350
rect 347278 28294 347334 28350
rect 347402 28294 347458 28350
rect 347526 28294 347582 28350
rect 347154 28170 347210 28226
rect 347278 28170 347334 28226
rect 347402 28170 347458 28226
rect 347526 28170 347582 28226
rect 347154 28046 347210 28102
rect 347278 28046 347334 28102
rect 347402 28046 347458 28102
rect 347526 28046 347582 28102
rect 347154 27922 347210 27978
rect 347278 27922 347334 27978
rect 347402 27922 347458 27978
rect 347526 27922 347582 27978
rect 347154 10294 347210 10350
rect 347278 10294 347334 10350
rect 347402 10294 347458 10350
rect 347526 10294 347582 10350
rect 347154 10170 347210 10226
rect 347278 10170 347334 10226
rect 347402 10170 347458 10226
rect 347526 10170 347582 10226
rect 347154 10046 347210 10102
rect 347278 10046 347334 10102
rect 347402 10046 347458 10102
rect 347526 10046 347582 10102
rect 347154 9922 347210 9978
rect 347278 9922 347334 9978
rect 347402 9922 347458 9978
rect 347526 9922 347582 9978
rect 350252 311642 350308 311698
rect 353612 324962 353668 325018
rect 374154 346294 374210 346350
rect 374278 346294 374334 346350
rect 374402 346294 374458 346350
rect 374526 346294 374582 346350
rect 374154 346170 374210 346226
rect 374278 346170 374334 346226
rect 374402 346170 374458 346226
rect 374526 346170 374582 346226
rect 374154 346046 374210 346102
rect 374278 346046 374334 346102
rect 374402 346046 374458 346102
rect 374526 346046 374582 346102
rect 374154 345922 374210 345978
rect 374278 345922 374334 345978
rect 374402 345922 374458 345978
rect 374526 345922 374582 345978
rect 358652 343682 358708 343738
rect 374154 328294 374210 328350
rect 374278 328294 374334 328350
rect 374402 328294 374458 328350
rect 374526 328294 374582 328350
rect 374154 328170 374210 328226
rect 374278 328170 374334 328226
rect 374402 328170 374458 328226
rect 374526 328170 374582 328226
rect 374154 328046 374210 328102
rect 374278 328046 374334 328102
rect 374402 328046 374458 328102
rect 374526 328046 374582 328102
rect 374154 327922 374210 327978
rect 374278 327922 374334 327978
rect 374402 327922 374458 327978
rect 374526 327922 374582 327978
rect 360332 323342 360388 323398
rect 374154 310294 374210 310350
rect 374278 310294 374334 310350
rect 374402 310294 374458 310350
rect 374526 310294 374582 310350
rect 374154 310170 374210 310226
rect 374278 310170 374334 310226
rect 374402 310170 374458 310226
rect 374526 310170 374582 310226
rect 374154 310046 374210 310102
rect 374278 310046 374334 310102
rect 374402 310046 374458 310102
rect 374526 310046 374582 310102
rect 374154 309922 374210 309978
rect 374278 309922 374334 309978
rect 374402 309922 374458 309978
rect 374526 309922 374582 309978
rect 374154 292294 374210 292350
rect 374278 292294 374334 292350
rect 374402 292294 374458 292350
rect 374526 292294 374582 292350
rect 374154 292170 374210 292226
rect 374278 292170 374334 292226
rect 374402 292170 374458 292226
rect 374526 292170 374582 292226
rect 374154 292046 374210 292102
rect 374278 292046 374334 292102
rect 374402 292046 374458 292102
rect 374526 292046 374582 292102
rect 374154 291922 374210 291978
rect 374278 291922 374334 291978
rect 374402 291922 374458 291978
rect 374526 291922 374582 291978
rect 374154 274294 374210 274350
rect 374278 274294 374334 274350
rect 374402 274294 374458 274350
rect 374526 274294 374582 274350
rect 374154 274170 374210 274226
rect 374278 274170 374334 274226
rect 374402 274170 374458 274226
rect 374526 274170 374582 274226
rect 374154 274046 374210 274102
rect 374278 274046 374334 274102
rect 374402 274046 374458 274102
rect 374526 274046 374582 274102
rect 374154 273922 374210 273978
rect 374278 273922 374334 273978
rect 374402 273922 374458 273978
rect 374526 273922 374582 273978
rect 361930 244294 361986 244350
rect 362054 244294 362110 244350
rect 362178 244294 362234 244350
rect 362302 244294 362358 244350
rect 361930 244170 361986 244226
rect 362054 244170 362110 244226
rect 362178 244170 362234 244226
rect 362302 244170 362358 244226
rect 361930 244046 361986 244102
rect 362054 244046 362110 244102
rect 362178 244046 362234 244102
rect 362302 244046 362358 244102
rect 361930 243922 361986 243978
rect 362054 243922 362110 243978
rect 362178 243922 362234 243978
rect 362302 243922 362358 243978
rect 361130 238294 361186 238350
rect 361254 238294 361310 238350
rect 361378 238294 361434 238350
rect 361502 238294 361558 238350
rect 361130 238170 361186 238226
rect 361254 238170 361310 238226
rect 361378 238170 361434 238226
rect 361502 238170 361558 238226
rect 361130 238046 361186 238102
rect 361254 238046 361310 238102
rect 361378 238046 361434 238102
rect 361502 238046 361558 238102
rect 361130 237922 361186 237978
rect 361254 237922 361310 237978
rect 361378 237922 361434 237978
rect 361502 237922 361558 237978
rect 361930 226294 361986 226350
rect 362054 226294 362110 226350
rect 362178 226294 362234 226350
rect 362302 226294 362358 226350
rect 361930 226170 361986 226226
rect 362054 226170 362110 226226
rect 362178 226170 362234 226226
rect 362302 226170 362358 226226
rect 361930 226046 361986 226102
rect 362054 226046 362110 226102
rect 362178 226046 362234 226102
rect 362302 226046 362358 226102
rect 361930 225922 361986 225978
rect 362054 225922 362110 225978
rect 362178 225922 362234 225978
rect 362302 225922 362358 225978
rect 361130 220294 361186 220350
rect 361254 220294 361310 220350
rect 361378 220294 361434 220350
rect 361502 220294 361558 220350
rect 361130 220170 361186 220226
rect 361254 220170 361310 220226
rect 361378 220170 361434 220226
rect 361502 220170 361558 220226
rect 361130 220046 361186 220102
rect 361254 220046 361310 220102
rect 361378 220046 361434 220102
rect 361502 220046 361558 220102
rect 361130 219922 361186 219978
rect 361254 219922 361310 219978
rect 361378 219922 361434 219978
rect 361502 219922 361558 219978
rect 361930 208294 361986 208350
rect 362054 208294 362110 208350
rect 362178 208294 362234 208350
rect 362302 208294 362358 208350
rect 361930 208170 361986 208226
rect 362054 208170 362110 208226
rect 362178 208170 362234 208226
rect 362302 208170 362358 208226
rect 361930 208046 361986 208102
rect 362054 208046 362110 208102
rect 362178 208046 362234 208102
rect 362302 208046 362358 208102
rect 361930 207922 361986 207978
rect 362054 207922 362110 207978
rect 362178 207922 362234 207978
rect 362302 207922 362358 207978
rect 361130 202294 361186 202350
rect 361254 202294 361310 202350
rect 361378 202294 361434 202350
rect 361502 202294 361558 202350
rect 361130 202170 361186 202226
rect 361254 202170 361310 202226
rect 361378 202170 361434 202226
rect 361502 202170 361558 202226
rect 361130 202046 361186 202102
rect 361254 202046 361310 202102
rect 361378 202046 361434 202102
rect 361502 202046 361558 202102
rect 361130 201922 361186 201978
rect 361254 201922 361310 201978
rect 361378 201922 361434 201978
rect 361502 201922 361558 201978
rect 361930 190294 361986 190350
rect 362054 190294 362110 190350
rect 362178 190294 362234 190350
rect 362302 190294 362358 190350
rect 361930 190170 361986 190226
rect 362054 190170 362110 190226
rect 362178 190170 362234 190226
rect 362302 190170 362358 190226
rect 361930 190046 361986 190102
rect 362054 190046 362110 190102
rect 362178 190046 362234 190102
rect 362302 190046 362358 190102
rect 361930 189922 361986 189978
rect 362054 189922 362110 189978
rect 362178 189922 362234 189978
rect 362302 189922 362358 189978
rect 361130 184294 361186 184350
rect 361254 184294 361310 184350
rect 361378 184294 361434 184350
rect 361502 184294 361558 184350
rect 361130 184170 361186 184226
rect 361254 184170 361310 184226
rect 361378 184170 361434 184226
rect 361502 184170 361558 184226
rect 361130 184046 361186 184102
rect 361254 184046 361310 184102
rect 361378 184046 361434 184102
rect 361502 184046 361558 184102
rect 361130 183922 361186 183978
rect 361254 183922 361310 183978
rect 361378 183922 361434 183978
rect 361502 183922 361558 183978
rect 361930 172294 361986 172350
rect 362054 172294 362110 172350
rect 362178 172294 362234 172350
rect 362302 172294 362358 172350
rect 361930 172170 361986 172226
rect 362054 172170 362110 172226
rect 362178 172170 362234 172226
rect 362302 172170 362358 172226
rect 361930 172046 361986 172102
rect 362054 172046 362110 172102
rect 362178 172046 362234 172102
rect 362302 172046 362358 172102
rect 361930 171922 361986 171978
rect 362054 171922 362110 171978
rect 362178 171922 362234 171978
rect 362302 171922 362358 171978
rect 361130 166294 361186 166350
rect 361254 166294 361310 166350
rect 361378 166294 361434 166350
rect 361502 166294 361558 166350
rect 361130 166170 361186 166226
rect 361254 166170 361310 166226
rect 361378 166170 361434 166226
rect 361502 166170 361558 166226
rect 361130 166046 361186 166102
rect 361254 166046 361310 166102
rect 361378 166046 361434 166102
rect 361502 166046 361558 166102
rect 361130 165922 361186 165978
rect 361254 165922 361310 165978
rect 361378 165922 361434 165978
rect 361502 165922 361558 165978
rect 377874 388294 377930 388350
rect 377998 388294 378054 388350
rect 378122 388294 378178 388350
rect 378246 388294 378302 388350
rect 377874 388170 377930 388226
rect 377998 388170 378054 388226
rect 378122 388170 378178 388226
rect 378246 388170 378302 388226
rect 377874 388046 377930 388102
rect 377998 388046 378054 388102
rect 378122 388046 378178 388102
rect 378246 388046 378302 388102
rect 377874 387922 377930 387978
rect 377998 387922 378054 387978
rect 378122 387922 378178 387978
rect 378246 387922 378302 387978
rect 404874 400294 404930 400350
rect 404998 400294 405054 400350
rect 405122 400294 405178 400350
rect 405246 400294 405302 400350
rect 404874 400170 404930 400226
rect 404998 400170 405054 400226
rect 405122 400170 405178 400226
rect 405246 400170 405302 400226
rect 404874 400046 404930 400102
rect 404998 400046 405054 400102
rect 405122 400046 405178 400102
rect 405246 400046 405302 400102
rect 404874 399922 404930 399978
rect 404998 399922 405054 399978
rect 405122 399922 405178 399978
rect 405246 399922 405302 399978
rect 404874 382294 404930 382350
rect 404998 382294 405054 382350
rect 405122 382294 405178 382350
rect 405246 382294 405302 382350
rect 404874 382170 404930 382226
rect 404998 382170 405054 382226
rect 405122 382170 405178 382226
rect 405246 382170 405302 382226
rect 404874 382046 404930 382102
rect 404998 382046 405054 382102
rect 405122 382046 405178 382102
rect 405246 382046 405302 382102
rect 404874 381922 404930 381978
rect 404998 381922 405054 381978
rect 405122 381922 405178 381978
rect 405246 381922 405302 381978
rect 377874 370294 377930 370350
rect 377998 370294 378054 370350
rect 378122 370294 378178 370350
rect 378246 370294 378302 370350
rect 377874 370170 377930 370226
rect 377998 370170 378054 370226
rect 378122 370170 378178 370226
rect 378246 370170 378302 370226
rect 377874 370046 377930 370102
rect 377998 370046 378054 370102
rect 378122 370046 378178 370102
rect 378246 370046 378302 370102
rect 377874 369922 377930 369978
rect 377998 369922 378054 369978
rect 378122 369922 378178 369978
rect 378246 369922 378302 369978
rect 386614 370294 386670 370350
rect 386738 370294 386794 370350
rect 386862 370294 386918 370350
rect 386986 370294 387042 370350
rect 386614 370170 386670 370226
rect 386738 370170 386794 370226
rect 386862 370170 386918 370226
rect 386986 370170 387042 370226
rect 386614 370046 386670 370102
rect 386738 370046 386794 370102
rect 386862 370046 386918 370102
rect 386986 370046 387042 370102
rect 386614 369922 386670 369978
rect 386738 369922 386794 369978
rect 386862 369922 386918 369978
rect 386986 369922 387042 369978
rect 387414 364294 387470 364350
rect 387538 364294 387594 364350
rect 387662 364294 387718 364350
rect 387786 364294 387842 364350
rect 387414 364170 387470 364226
rect 387538 364170 387594 364226
rect 387662 364170 387718 364226
rect 387786 364170 387842 364226
rect 387414 364046 387470 364102
rect 387538 364046 387594 364102
rect 387662 364046 387718 364102
rect 387786 364046 387842 364102
rect 387414 363922 387470 363978
rect 387538 363922 387594 363978
rect 387662 363922 387718 363978
rect 387786 363922 387842 363978
rect 404874 364294 404930 364350
rect 404998 364294 405054 364350
rect 405122 364294 405178 364350
rect 405246 364294 405302 364350
rect 404874 364170 404930 364226
rect 404998 364170 405054 364226
rect 405122 364170 405178 364226
rect 405246 364170 405302 364226
rect 404874 364046 404930 364102
rect 404998 364046 405054 364102
rect 405122 364046 405178 364102
rect 405246 364046 405302 364102
rect 404874 363922 404930 363978
rect 404998 363922 405054 363978
rect 405122 363922 405178 363978
rect 405246 363922 405302 363978
rect 377874 352294 377930 352350
rect 377998 352294 378054 352350
rect 378122 352294 378178 352350
rect 378246 352294 378302 352350
rect 377874 352170 377930 352226
rect 377998 352170 378054 352226
rect 378122 352170 378178 352226
rect 378246 352170 378302 352226
rect 377874 352046 377930 352102
rect 377998 352046 378054 352102
rect 378122 352046 378178 352102
rect 378246 352046 378302 352102
rect 377874 351922 377930 351978
rect 377998 351922 378054 351978
rect 378122 351922 378178 351978
rect 378246 351922 378302 351978
rect 386614 352294 386670 352350
rect 386738 352294 386794 352350
rect 386862 352294 386918 352350
rect 386986 352294 387042 352350
rect 386614 352170 386670 352226
rect 386738 352170 386794 352226
rect 386862 352170 386918 352226
rect 386986 352170 387042 352226
rect 386614 352046 386670 352102
rect 386738 352046 386794 352102
rect 386862 352046 386918 352102
rect 386986 352046 387042 352102
rect 386614 351922 386670 351978
rect 386738 351922 386794 351978
rect 386862 351922 386918 351978
rect 386986 351922 387042 351978
rect 387414 346294 387470 346350
rect 387538 346294 387594 346350
rect 387662 346294 387718 346350
rect 387786 346294 387842 346350
rect 387414 346170 387470 346226
rect 387538 346170 387594 346226
rect 387662 346170 387718 346226
rect 387786 346170 387842 346226
rect 387414 346046 387470 346102
rect 387538 346046 387594 346102
rect 387662 346046 387718 346102
rect 387786 346046 387842 346102
rect 387414 345922 387470 345978
rect 387538 345922 387594 345978
rect 387662 345922 387718 345978
rect 387786 345922 387842 345978
rect 404874 346294 404930 346350
rect 404998 346294 405054 346350
rect 405122 346294 405178 346350
rect 405246 346294 405302 346350
rect 404874 346170 404930 346226
rect 404998 346170 405054 346226
rect 405122 346170 405178 346226
rect 405246 346170 405302 346226
rect 404874 346046 404930 346102
rect 404998 346046 405054 346102
rect 405122 346046 405178 346102
rect 405246 346046 405302 346102
rect 404874 345922 404930 345978
rect 404998 345922 405054 345978
rect 405122 345922 405178 345978
rect 405246 345922 405302 345978
rect 377874 334294 377930 334350
rect 377998 334294 378054 334350
rect 378122 334294 378178 334350
rect 378246 334294 378302 334350
rect 377874 334170 377930 334226
rect 377998 334170 378054 334226
rect 378122 334170 378178 334226
rect 378246 334170 378302 334226
rect 377874 334046 377930 334102
rect 377998 334046 378054 334102
rect 378122 334046 378178 334102
rect 378246 334046 378302 334102
rect 377874 333922 377930 333978
rect 377998 333922 378054 333978
rect 378122 333922 378178 333978
rect 378246 333922 378302 333978
rect 386614 334294 386670 334350
rect 386738 334294 386794 334350
rect 386862 334294 386918 334350
rect 386986 334294 387042 334350
rect 386614 334170 386670 334226
rect 386738 334170 386794 334226
rect 386862 334170 386918 334226
rect 386986 334170 387042 334226
rect 386614 334046 386670 334102
rect 386738 334046 386794 334102
rect 386862 334046 386918 334102
rect 386986 334046 387042 334102
rect 386614 333922 386670 333978
rect 386738 333922 386794 333978
rect 386862 333922 386918 333978
rect 386986 333922 387042 333978
rect 387414 328294 387470 328350
rect 387538 328294 387594 328350
rect 387662 328294 387718 328350
rect 387786 328294 387842 328350
rect 387414 328170 387470 328226
rect 387538 328170 387594 328226
rect 387662 328170 387718 328226
rect 387786 328170 387842 328226
rect 387414 328046 387470 328102
rect 387538 328046 387594 328102
rect 387662 328046 387718 328102
rect 387786 328046 387842 328102
rect 387414 327922 387470 327978
rect 387538 327922 387594 327978
rect 387662 327922 387718 327978
rect 387786 327922 387842 327978
rect 377874 316294 377930 316350
rect 377998 316294 378054 316350
rect 378122 316294 378178 316350
rect 378246 316294 378302 316350
rect 377874 316170 377930 316226
rect 377998 316170 378054 316226
rect 378122 316170 378178 316226
rect 378246 316170 378302 316226
rect 377874 316046 377930 316102
rect 377998 316046 378054 316102
rect 378122 316046 378178 316102
rect 378246 316046 378302 316102
rect 377874 315922 377930 315978
rect 377998 315922 378054 315978
rect 378122 315922 378178 315978
rect 378246 315922 378302 315978
rect 386614 316294 386670 316350
rect 386738 316294 386794 316350
rect 386862 316294 386918 316350
rect 386986 316294 387042 316350
rect 386614 316170 386670 316226
rect 386738 316170 386794 316226
rect 386862 316170 386918 316226
rect 386986 316170 387042 316226
rect 386614 316046 386670 316102
rect 386738 316046 386794 316102
rect 386862 316046 386918 316102
rect 386986 316046 387042 316102
rect 386614 315922 386670 315978
rect 386738 315922 386794 315978
rect 386862 315922 386918 315978
rect 386986 315922 387042 315978
rect 387414 310294 387470 310350
rect 387538 310294 387594 310350
rect 387662 310294 387718 310350
rect 387786 310294 387842 310350
rect 387414 310170 387470 310226
rect 387538 310170 387594 310226
rect 387662 310170 387718 310226
rect 387786 310170 387842 310226
rect 387414 310046 387470 310102
rect 387538 310046 387594 310102
rect 387662 310046 387718 310102
rect 387786 310046 387842 310102
rect 387414 309922 387470 309978
rect 387538 309922 387594 309978
rect 387662 309922 387718 309978
rect 387786 309922 387842 309978
rect 387996 301742 388052 301798
rect 387996 300302 388052 300358
rect 388220 300302 388276 300358
rect 377874 298294 377930 298350
rect 377998 298294 378054 298350
rect 378122 298294 378178 298350
rect 378246 298294 378302 298350
rect 377874 298170 377930 298226
rect 377998 298170 378054 298226
rect 378122 298170 378178 298226
rect 378246 298170 378302 298226
rect 377874 298046 377930 298102
rect 377998 298046 378054 298102
rect 378122 298046 378178 298102
rect 378246 298046 378302 298102
rect 377874 297922 377930 297978
rect 377998 297922 378054 297978
rect 378122 297922 378178 297978
rect 378246 297922 378302 297978
rect 386614 298294 386670 298350
rect 386738 298294 386794 298350
rect 386862 298294 386918 298350
rect 386986 298294 387042 298350
rect 386614 298170 386670 298226
rect 386738 298170 386794 298226
rect 386862 298170 386918 298226
rect 386986 298170 387042 298226
rect 386614 298046 386670 298102
rect 386738 298046 386794 298102
rect 386862 298046 386918 298102
rect 386986 298046 387042 298102
rect 386614 297922 386670 297978
rect 386738 297922 386794 297978
rect 386862 297922 386918 297978
rect 386986 297922 387042 297978
rect 390572 297062 390628 297118
rect 404874 328294 404930 328350
rect 404998 328294 405054 328350
rect 405122 328294 405178 328350
rect 405246 328294 405302 328350
rect 404874 328170 404930 328226
rect 404998 328170 405054 328226
rect 405122 328170 405178 328226
rect 405246 328170 405302 328226
rect 404874 328046 404930 328102
rect 404998 328046 405054 328102
rect 405122 328046 405178 328102
rect 405246 328046 405302 328102
rect 404874 327922 404930 327978
rect 404998 327922 405054 327978
rect 405122 327922 405178 327978
rect 405246 327922 405302 327978
rect 404874 310294 404930 310350
rect 404998 310294 405054 310350
rect 405122 310294 405178 310350
rect 405246 310294 405302 310350
rect 404874 310170 404930 310226
rect 404998 310170 405054 310226
rect 405122 310170 405178 310226
rect 405246 310170 405302 310226
rect 404874 310046 404930 310102
rect 404998 310046 405054 310102
rect 405122 310046 405178 310102
rect 405246 310046 405302 310102
rect 404874 309922 404930 309978
rect 404998 309922 405054 309978
rect 405122 309922 405178 309978
rect 405246 309922 405302 309978
rect 388444 296882 388500 296938
rect 387996 296702 388052 296758
rect 387414 292294 387470 292350
rect 387538 292294 387594 292350
rect 387662 292294 387718 292350
rect 387786 292294 387842 292350
rect 387414 292170 387470 292226
rect 387538 292170 387594 292226
rect 387662 292170 387718 292226
rect 387786 292170 387842 292226
rect 387414 292046 387470 292102
rect 387538 292046 387594 292102
rect 387662 292046 387718 292102
rect 387786 292046 387842 292102
rect 387414 291922 387470 291978
rect 387538 291922 387594 291978
rect 387662 291922 387718 291978
rect 387786 291922 387842 291978
rect 404874 292294 404930 292350
rect 404998 292294 405054 292350
rect 405122 292294 405178 292350
rect 405246 292294 405302 292350
rect 387996 291662 388052 291718
rect 404874 292170 404930 292226
rect 404998 292170 405054 292226
rect 405122 292170 405178 292226
rect 405246 292170 405302 292226
rect 404874 292046 404930 292102
rect 404998 292046 405054 292102
rect 405122 292046 405178 292102
rect 405246 292046 405302 292102
rect 404874 291922 404930 291978
rect 404998 291922 405054 291978
rect 405122 291922 405178 291978
rect 405246 291922 405302 291978
rect 387996 290222 388052 290278
rect 377874 280294 377930 280350
rect 377998 280294 378054 280350
rect 378122 280294 378178 280350
rect 378246 280294 378302 280350
rect 377874 280170 377930 280226
rect 377998 280170 378054 280226
rect 378122 280170 378178 280226
rect 378246 280170 378302 280226
rect 377874 280046 377930 280102
rect 377998 280046 378054 280102
rect 378122 280046 378178 280102
rect 378246 280046 378302 280102
rect 377874 279922 377930 279978
rect 377998 279922 378054 279978
rect 378122 279922 378178 279978
rect 378246 279922 378302 279978
rect 377874 262294 377930 262350
rect 377998 262294 378054 262350
rect 378122 262294 378178 262350
rect 378246 262294 378302 262350
rect 377874 262170 377930 262226
rect 377998 262170 378054 262226
rect 378122 262170 378178 262226
rect 378246 262170 378302 262226
rect 377874 262046 377930 262102
rect 377998 262046 378054 262102
rect 378122 262046 378178 262102
rect 378246 262046 378302 262102
rect 377874 261922 377930 261978
rect 377998 261922 378054 261978
rect 378122 261922 378178 261978
rect 378246 261922 378302 261978
rect 374154 256294 374210 256350
rect 374278 256294 374334 256350
rect 374402 256294 374458 256350
rect 374526 256294 374582 256350
rect 374154 256170 374210 256226
rect 374278 256170 374334 256226
rect 374402 256170 374458 256226
rect 374526 256170 374582 256226
rect 374154 256046 374210 256102
rect 374278 256046 374334 256102
rect 374402 256046 374458 256102
rect 374526 256046 374582 256102
rect 374154 255922 374210 255978
rect 374278 255922 374334 255978
rect 374402 255922 374458 255978
rect 374526 255922 374582 255978
rect 374154 238294 374210 238350
rect 374278 238294 374334 238350
rect 374402 238294 374458 238350
rect 374526 238294 374582 238350
rect 374154 238170 374210 238226
rect 374278 238170 374334 238226
rect 374402 238170 374458 238226
rect 374526 238170 374582 238226
rect 374154 238046 374210 238102
rect 374278 238046 374334 238102
rect 374402 238046 374458 238102
rect 374526 238046 374582 238102
rect 374154 237922 374210 237978
rect 374278 237922 374334 237978
rect 374402 237922 374458 237978
rect 374526 237922 374582 237978
rect 374154 220294 374210 220350
rect 374278 220294 374334 220350
rect 374402 220294 374458 220350
rect 374526 220294 374582 220350
rect 374154 220170 374210 220226
rect 374278 220170 374334 220226
rect 374402 220170 374458 220226
rect 374526 220170 374582 220226
rect 374154 220046 374210 220102
rect 374278 220046 374334 220102
rect 374402 220046 374458 220102
rect 374526 220046 374582 220102
rect 374154 219922 374210 219978
rect 374278 219922 374334 219978
rect 374402 219922 374458 219978
rect 374526 219922 374582 219978
rect 374154 202294 374210 202350
rect 374278 202294 374334 202350
rect 374402 202294 374458 202350
rect 374526 202294 374582 202350
rect 374154 202170 374210 202226
rect 374278 202170 374334 202226
rect 374402 202170 374458 202226
rect 374526 202170 374582 202226
rect 374154 202046 374210 202102
rect 374278 202046 374334 202102
rect 374402 202046 374458 202102
rect 374526 202046 374582 202102
rect 374154 201922 374210 201978
rect 374278 201922 374334 201978
rect 374402 201922 374458 201978
rect 374526 201922 374582 201978
rect 374154 184294 374210 184350
rect 374278 184294 374334 184350
rect 374402 184294 374458 184350
rect 374526 184294 374582 184350
rect 374154 184170 374210 184226
rect 374278 184170 374334 184226
rect 374402 184170 374458 184226
rect 374526 184170 374582 184226
rect 374154 184046 374210 184102
rect 374278 184046 374334 184102
rect 374402 184046 374458 184102
rect 374526 184046 374582 184102
rect 374154 183922 374210 183978
rect 374278 183922 374334 183978
rect 374402 183922 374458 183978
rect 374526 183922 374582 183978
rect 374154 166294 374210 166350
rect 374278 166294 374334 166350
rect 374402 166294 374458 166350
rect 374526 166294 374582 166350
rect 374154 166170 374210 166226
rect 374278 166170 374334 166226
rect 374402 166170 374458 166226
rect 374526 166170 374582 166226
rect 374154 166046 374210 166102
rect 374278 166046 374334 166102
rect 374402 166046 374458 166102
rect 374526 166046 374582 166102
rect 374154 165922 374210 165978
rect 374278 165922 374334 165978
rect 374402 165922 374458 165978
rect 374526 165922 374582 165978
rect 374154 148294 374210 148350
rect 374278 148294 374334 148350
rect 374402 148294 374458 148350
rect 374526 148294 374582 148350
rect 374154 148170 374210 148226
rect 374278 148170 374334 148226
rect 374402 148170 374458 148226
rect 374526 148170 374582 148226
rect 374154 148046 374210 148102
rect 374278 148046 374334 148102
rect 374402 148046 374458 148102
rect 374526 148046 374582 148102
rect 374154 147922 374210 147978
rect 374278 147922 374334 147978
rect 374402 147922 374458 147978
rect 374526 147922 374582 147978
rect 361130 130294 361186 130350
rect 361254 130294 361310 130350
rect 361378 130294 361434 130350
rect 361502 130294 361558 130350
rect 361130 130170 361186 130226
rect 361254 130170 361310 130226
rect 361378 130170 361434 130226
rect 361502 130170 361558 130226
rect 361130 130046 361186 130102
rect 361254 130046 361310 130102
rect 361378 130046 361434 130102
rect 361502 130046 361558 130102
rect 361130 129922 361186 129978
rect 361254 129922 361310 129978
rect 361378 129922 361434 129978
rect 361502 129922 361558 129978
rect 404874 274294 404930 274350
rect 404998 274294 405054 274350
rect 405122 274294 405178 274350
rect 405246 274294 405302 274350
rect 404874 274170 404930 274226
rect 404998 274170 405054 274226
rect 405122 274170 405178 274226
rect 405246 274170 405302 274226
rect 404874 274046 404930 274102
rect 404998 274046 405054 274102
rect 405122 274046 405178 274102
rect 405246 274046 405302 274102
rect 404874 273922 404930 273978
rect 404998 273922 405054 273978
rect 405122 273922 405178 273978
rect 405246 273922 405302 273978
rect 377874 244294 377930 244350
rect 377998 244294 378054 244350
rect 378122 244294 378178 244350
rect 378246 244294 378302 244350
rect 377874 244170 377930 244226
rect 377998 244170 378054 244226
rect 378122 244170 378178 244226
rect 378246 244170 378302 244226
rect 377874 244046 377930 244102
rect 377998 244046 378054 244102
rect 378122 244046 378178 244102
rect 378246 244046 378302 244102
rect 377874 243922 377930 243978
rect 377998 243922 378054 243978
rect 378122 243922 378178 243978
rect 378246 243922 378302 243978
rect 377874 226294 377930 226350
rect 377998 226294 378054 226350
rect 378122 226294 378178 226350
rect 378246 226294 378302 226350
rect 377874 226170 377930 226226
rect 377998 226170 378054 226226
rect 378122 226170 378178 226226
rect 378246 226170 378302 226226
rect 377874 226046 377930 226102
rect 377998 226046 378054 226102
rect 378122 226046 378178 226102
rect 378246 226046 378302 226102
rect 377874 225922 377930 225978
rect 377998 225922 378054 225978
rect 378122 225922 378178 225978
rect 378246 225922 378302 225978
rect 377874 208294 377930 208350
rect 377998 208294 378054 208350
rect 378122 208294 378178 208350
rect 378246 208294 378302 208350
rect 377874 208170 377930 208226
rect 377998 208170 378054 208226
rect 378122 208170 378178 208226
rect 378246 208170 378302 208226
rect 377874 208046 377930 208102
rect 377998 208046 378054 208102
rect 378122 208046 378178 208102
rect 378246 208046 378302 208102
rect 377874 207922 377930 207978
rect 377998 207922 378054 207978
rect 378122 207922 378178 207978
rect 378246 207922 378302 207978
rect 377874 190294 377930 190350
rect 377998 190294 378054 190350
rect 378122 190294 378178 190350
rect 378246 190294 378302 190350
rect 377874 190170 377930 190226
rect 377998 190170 378054 190226
rect 378122 190170 378178 190226
rect 378246 190170 378302 190226
rect 377874 190046 377930 190102
rect 377998 190046 378054 190102
rect 378122 190046 378178 190102
rect 378246 190046 378302 190102
rect 377874 189922 377930 189978
rect 377998 189922 378054 189978
rect 378122 189922 378178 189978
rect 378246 189922 378302 189978
rect 377874 172294 377930 172350
rect 377998 172294 378054 172350
rect 378122 172294 378178 172350
rect 378246 172294 378302 172350
rect 377874 172170 377930 172226
rect 377998 172170 378054 172226
rect 378122 172170 378178 172226
rect 378246 172170 378302 172226
rect 377874 172046 377930 172102
rect 377998 172046 378054 172102
rect 378122 172046 378178 172102
rect 378246 172046 378302 172102
rect 377874 171922 377930 171978
rect 377998 171922 378054 171978
rect 378122 171922 378178 171978
rect 378246 171922 378302 171978
rect 377874 154294 377930 154350
rect 377998 154294 378054 154350
rect 378122 154294 378178 154350
rect 378246 154294 378302 154350
rect 377874 154170 377930 154226
rect 377998 154170 378054 154226
rect 378122 154170 378178 154226
rect 378246 154170 378302 154226
rect 377874 154046 377930 154102
rect 377998 154046 378054 154102
rect 378122 154046 378178 154102
rect 378246 154046 378302 154102
rect 377874 153922 377930 153978
rect 377998 153922 378054 153978
rect 378122 153922 378178 153978
rect 378246 153922 378302 153978
rect 374154 130294 374210 130350
rect 374278 130294 374334 130350
rect 374402 130294 374458 130350
rect 374526 130294 374582 130350
rect 374154 130170 374210 130226
rect 374278 130170 374334 130226
rect 374402 130170 374458 130226
rect 374526 130170 374582 130226
rect 374154 130046 374210 130102
rect 374278 130046 374334 130102
rect 374402 130046 374458 130102
rect 374526 130046 374582 130102
rect 374154 129922 374210 129978
rect 374278 129922 374334 129978
rect 374402 129922 374458 129978
rect 374526 129922 374582 129978
rect 361930 118294 361986 118350
rect 362054 118294 362110 118350
rect 362178 118294 362234 118350
rect 362302 118294 362358 118350
rect 361930 118170 361986 118226
rect 362054 118170 362110 118226
rect 362178 118170 362234 118226
rect 362302 118170 362358 118226
rect 361930 118046 361986 118102
rect 362054 118046 362110 118102
rect 362178 118046 362234 118102
rect 362302 118046 362358 118102
rect 361930 117922 361986 117978
rect 362054 117922 362110 117978
rect 362178 117922 362234 117978
rect 362302 117922 362358 117978
rect 361130 112294 361186 112350
rect 361254 112294 361310 112350
rect 361378 112294 361434 112350
rect 361502 112294 361558 112350
rect 361130 112170 361186 112226
rect 361254 112170 361310 112226
rect 361378 112170 361434 112226
rect 361502 112170 361558 112226
rect 361130 112046 361186 112102
rect 361254 112046 361310 112102
rect 361378 112046 361434 112102
rect 361502 112046 361558 112102
rect 361130 111922 361186 111978
rect 361254 111922 361310 111978
rect 361378 111922 361434 111978
rect 361502 111922 361558 111978
rect 374154 112294 374210 112350
rect 374278 112294 374334 112350
rect 374402 112294 374458 112350
rect 374526 112294 374582 112350
rect 374154 112170 374210 112226
rect 374278 112170 374334 112226
rect 374402 112170 374458 112226
rect 374526 112170 374582 112226
rect 374154 112046 374210 112102
rect 374278 112046 374334 112102
rect 374402 112046 374458 112102
rect 374526 112046 374582 112102
rect 374154 111922 374210 111978
rect 374278 111922 374334 111978
rect 374402 111922 374458 111978
rect 374526 111922 374582 111978
rect 361930 100294 361986 100350
rect 362054 100294 362110 100350
rect 362178 100294 362234 100350
rect 362302 100294 362358 100350
rect 361930 100170 361986 100226
rect 362054 100170 362110 100226
rect 362178 100170 362234 100226
rect 362302 100170 362358 100226
rect 361930 100046 361986 100102
rect 362054 100046 362110 100102
rect 362178 100046 362234 100102
rect 362302 100046 362358 100102
rect 361930 99922 361986 99978
rect 362054 99922 362110 99978
rect 362178 99922 362234 99978
rect 362302 99922 362358 99978
rect 361130 94294 361186 94350
rect 361254 94294 361310 94350
rect 361378 94294 361434 94350
rect 361502 94294 361558 94350
rect 361130 94170 361186 94226
rect 361254 94170 361310 94226
rect 361378 94170 361434 94226
rect 361502 94170 361558 94226
rect 361130 94046 361186 94102
rect 361254 94046 361310 94102
rect 361378 94046 361434 94102
rect 361502 94046 361558 94102
rect 361130 93922 361186 93978
rect 361254 93922 361310 93978
rect 361378 93922 361434 93978
rect 361502 93922 361558 93978
rect 374154 94294 374210 94350
rect 374278 94294 374334 94350
rect 374402 94294 374458 94350
rect 374526 94294 374582 94350
rect 374154 94170 374210 94226
rect 374278 94170 374334 94226
rect 374402 94170 374458 94226
rect 374526 94170 374582 94226
rect 374154 94046 374210 94102
rect 374278 94046 374334 94102
rect 374402 94046 374458 94102
rect 374526 94046 374582 94102
rect 374154 93922 374210 93978
rect 374278 93922 374334 93978
rect 374402 93922 374458 93978
rect 374526 93922 374582 93978
rect 361930 82294 361986 82350
rect 362054 82294 362110 82350
rect 362178 82294 362234 82350
rect 362302 82294 362358 82350
rect 361930 82170 361986 82226
rect 362054 82170 362110 82226
rect 362178 82170 362234 82226
rect 362302 82170 362358 82226
rect 361930 82046 361986 82102
rect 362054 82046 362110 82102
rect 362178 82046 362234 82102
rect 362302 82046 362358 82102
rect 361930 81922 361986 81978
rect 362054 81922 362110 81978
rect 362178 81922 362234 81978
rect 362302 81922 362358 81978
rect 361130 76294 361186 76350
rect 361254 76294 361310 76350
rect 361378 76294 361434 76350
rect 361502 76294 361558 76350
rect 361130 76170 361186 76226
rect 361254 76170 361310 76226
rect 361378 76170 361434 76226
rect 361502 76170 361558 76226
rect 361130 76046 361186 76102
rect 361254 76046 361310 76102
rect 361378 76046 361434 76102
rect 361502 76046 361558 76102
rect 361130 75922 361186 75978
rect 361254 75922 361310 75978
rect 361378 75922 361434 75978
rect 361502 75922 361558 75978
rect 374154 76294 374210 76350
rect 374278 76294 374334 76350
rect 374402 76294 374458 76350
rect 374526 76294 374582 76350
rect 374154 76170 374210 76226
rect 374278 76170 374334 76226
rect 374402 76170 374458 76226
rect 374526 76170 374582 76226
rect 374154 76046 374210 76102
rect 374278 76046 374334 76102
rect 374402 76046 374458 76102
rect 374526 76046 374582 76102
rect 374154 75922 374210 75978
rect 374278 75922 374334 75978
rect 374402 75922 374458 75978
rect 374526 75922 374582 75978
rect 361930 64294 361986 64350
rect 362054 64294 362110 64350
rect 362178 64294 362234 64350
rect 362302 64294 362358 64350
rect 361930 64170 361986 64226
rect 362054 64170 362110 64226
rect 362178 64170 362234 64226
rect 362302 64170 362358 64226
rect 361930 64046 361986 64102
rect 362054 64046 362110 64102
rect 362178 64046 362234 64102
rect 362302 64046 362358 64102
rect 361930 63922 361986 63978
rect 362054 63922 362110 63978
rect 362178 63922 362234 63978
rect 362302 63922 362358 63978
rect 361130 58294 361186 58350
rect 361254 58294 361310 58350
rect 361378 58294 361434 58350
rect 361502 58294 361558 58350
rect 361130 58170 361186 58226
rect 361254 58170 361310 58226
rect 361378 58170 361434 58226
rect 361502 58170 361558 58226
rect 361130 58046 361186 58102
rect 361254 58046 361310 58102
rect 361378 58046 361434 58102
rect 361502 58046 361558 58102
rect 361130 57922 361186 57978
rect 361254 57922 361310 57978
rect 361378 57922 361434 57978
rect 361502 57922 361558 57978
rect 374154 58294 374210 58350
rect 374278 58294 374334 58350
rect 374402 58294 374458 58350
rect 374526 58294 374582 58350
rect 374154 58170 374210 58226
rect 374278 58170 374334 58226
rect 374402 58170 374458 58226
rect 374526 58170 374582 58226
rect 374154 58046 374210 58102
rect 374278 58046 374334 58102
rect 374402 58046 374458 58102
rect 374526 58046 374582 58102
rect 374154 57922 374210 57978
rect 374278 57922 374334 57978
rect 374402 57922 374458 57978
rect 374526 57922 374582 57978
rect 361930 46294 361986 46350
rect 362054 46294 362110 46350
rect 362178 46294 362234 46350
rect 362302 46294 362358 46350
rect 361930 46170 361986 46226
rect 362054 46170 362110 46226
rect 362178 46170 362234 46226
rect 362302 46170 362358 46226
rect 361930 46046 361986 46102
rect 362054 46046 362110 46102
rect 362178 46046 362234 46102
rect 362302 46046 362358 46102
rect 361930 45922 361986 45978
rect 362054 45922 362110 45978
rect 362178 45922 362234 45978
rect 362302 45922 362358 45978
rect 374154 40294 374210 40350
rect 374278 40294 374334 40350
rect 374402 40294 374458 40350
rect 374526 40294 374582 40350
rect 374154 40170 374210 40226
rect 374278 40170 374334 40226
rect 374402 40170 374458 40226
rect 374526 40170 374582 40226
rect 374154 40046 374210 40102
rect 374278 40046 374334 40102
rect 374402 40046 374458 40102
rect 374526 40046 374582 40102
rect 374154 39922 374210 39978
rect 374278 39922 374334 39978
rect 374402 39922 374458 39978
rect 374526 39922 374582 39978
rect 374154 22294 374210 22350
rect 374278 22294 374334 22350
rect 374402 22294 374458 22350
rect 374526 22294 374582 22350
rect 374154 22170 374210 22226
rect 374278 22170 374334 22226
rect 374402 22170 374458 22226
rect 374526 22170 374582 22226
rect 374154 22046 374210 22102
rect 374278 22046 374334 22102
rect 374402 22046 374458 22102
rect 374526 22046 374582 22102
rect 374154 21922 374210 21978
rect 374278 21922 374334 21978
rect 374402 21922 374458 21978
rect 374526 21922 374582 21978
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 347154 -1176 347210 -1120
rect 347278 -1176 347334 -1120
rect 347402 -1176 347458 -1120
rect 347526 -1176 347582 -1120
rect 347154 -1300 347210 -1244
rect 347278 -1300 347334 -1244
rect 347402 -1300 347458 -1244
rect 347526 -1300 347582 -1244
rect 347154 -1424 347210 -1368
rect 347278 -1424 347334 -1368
rect 347402 -1424 347458 -1368
rect 347526 -1424 347582 -1368
rect 347154 -1548 347210 -1492
rect 347278 -1548 347334 -1492
rect 347402 -1548 347458 -1492
rect 347526 -1548 347582 -1492
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 404874 256294 404930 256350
rect 404998 256294 405054 256350
rect 405122 256294 405178 256350
rect 405246 256294 405302 256350
rect 404874 256170 404930 256226
rect 404998 256170 405054 256226
rect 405122 256170 405178 256226
rect 405246 256170 405302 256226
rect 404874 256046 404930 256102
rect 404998 256046 405054 256102
rect 405122 256046 405178 256102
rect 405246 256046 405302 256102
rect 404874 255922 404930 255978
rect 404998 255922 405054 255978
rect 405122 255922 405178 255978
rect 405246 255922 405302 255978
rect 404874 238294 404930 238350
rect 404998 238294 405054 238350
rect 405122 238294 405178 238350
rect 405246 238294 405302 238350
rect 404874 238170 404930 238226
rect 404998 238170 405054 238226
rect 405122 238170 405178 238226
rect 405246 238170 405302 238226
rect 404874 238046 404930 238102
rect 404998 238046 405054 238102
rect 405122 238046 405178 238102
rect 405246 238046 405302 238102
rect 404874 237922 404930 237978
rect 404998 237922 405054 237978
rect 405122 237922 405178 237978
rect 405246 237922 405302 237978
rect 404874 220294 404930 220350
rect 404998 220294 405054 220350
rect 405122 220294 405178 220350
rect 405246 220294 405302 220350
rect 404874 220170 404930 220226
rect 404998 220170 405054 220226
rect 405122 220170 405178 220226
rect 405246 220170 405302 220226
rect 404874 220046 404930 220102
rect 404998 220046 405054 220102
rect 405122 220046 405178 220102
rect 405246 220046 405302 220102
rect 404874 219922 404930 219978
rect 404998 219922 405054 219978
rect 405122 219922 405178 219978
rect 405246 219922 405302 219978
rect 404874 202294 404930 202350
rect 404998 202294 405054 202350
rect 405122 202294 405178 202350
rect 405246 202294 405302 202350
rect 404874 202170 404930 202226
rect 404998 202170 405054 202226
rect 405122 202170 405178 202226
rect 405246 202170 405302 202226
rect 404874 202046 404930 202102
rect 404998 202046 405054 202102
rect 405122 202046 405178 202102
rect 405246 202046 405302 202102
rect 404874 201922 404930 201978
rect 404998 201922 405054 201978
rect 405122 201922 405178 201978
rect 405246 201922 405302 201978
rect 404874 184294 404930 184350
rect 404998 184294 405054 184350
rect 405122 184294 405178 184350
rect 405246 184294 405302 184350
rect 404874 184170 404930 184226
rect 404998 184170 405054 184226
rect 405122 184170 405178 184226
rect 405246 184170 405302 184226
rect 404874 184046 404930 184102
rect 404998 184046 405054 184102
rect 405122 184046 405178 184102
rect 405246 184046 405302 184102
rect 404874 183922 404930 183978
rect 404998 183922 405054 183978
rect 405122 183922 405178 183978
rect 405246 183922 405302 183978
rect 404874 166294 404930 166350
rect 404998 166294 405054 166350
rect 405122 166294 405178 166350
rect 405246 166294 405302 166350
rect 404874 166170 404930 166226
rect 404998 166170 405054 166226
rect 405122 166170 405178 166226
rect 405246 166170 405302 166226
rect 404874 166046 404930 166102
rect 404998 166046 405054 166102
rect 405122 166046 405178 166102
rect 405246 166046 405302 166102
rect 404874 165922 404930 165978
rect 404998 165922 405054 165978
rect 405122 165922 405178 165978
rect 405246 165922 405302 165978
rect 404874 148294 404930 148350
rect 404998 148294 405054 148350
rect 405122 148294 405178 148350
rect 405246 148294 405302 148350
rect 404874 148170 404930 148226
rect 404998 148170 405054 148226
rect 405122 148170 405178 148226
rect 405246 148170 405302 148226
rect 404874 148046 404930 148102
rect 404998 148046 405054 148102
rect 405122 148046 405178 148102
rect 405246 148046 405302 148102
rect 404874 147922 404930 147978
rect 404998 147922 405054 147978
rect 405122 147922 405178 147978
rect 405246 147922 405302 147978
rect 377874 136294 377930 136350
rect 377998 136294 378054 136350
rect 378122 136294 378178 136350
rect 378246 136294 378302 136350
rect 377874 136170 377930 136226
rect 377998 136170 378054 136226
rect 378122 136170 378178 136226
rect 378246 136170 378302 136226
rect 377874 136046 377930 136102
rect 377998 136046 378054 136102
rect 378122 136046 378178 136102
rect 378246 136046 378302 136102
rect 377874 135922 377930 135978
rect 377998 135922 378054 135978
rect 378122 135922 378178 135978
rect 378246 135922 378302 135978
rect 377874 118294 377930 118350
rect 377998 118294 378054 118350
rect 378122 118294 378178 118350
rect 378246 118294 378302 118350
rect 377874 118170 377930 118226
rect 377998 118170 378054 118226
rect 378122 118170 378178 118226
rect 378246 118170 378302 118226
rect 377874 118046 377930 118102
rect 377998 118046 378054 118102
rect 378122 118046 378178 118102
rect 378246 118046 378302 118102
rect 377874 117922 377930 117978
rect 377998 117922 378054 117978
rect 378122 117922 378178 117978
rect 378246 117922 378302 117978
rect 377874 100294 377930 100350
rect 377998 100294 378054 100350
rect 378122 100294 378178 100350
rect 378246 100294 378302 100350
rect 377874 100170 377930 100226
rect 377998 100170 378054 100226
rect 378122 100170 378178 100226
rect 378246 100170 378302 100226
rect 377874 100046 377930 100102
rect 377998 100046 378054 100102
rect 378122 100046 378178 100102
rect 378246 100046 378302 100102
rect 377874 99922 377930 99978
rect 377998 99922 378054 99978
rect 378122 99922 378178 99978
rect 378246 99922 378302 99978
rect 377874 82294 377930 82350
rect 377998 82294 378054 82350
rect 378122 82294 378178 82350
rect 378246 82294 378302 82350
rect 377874 82170 377930 82226
rect 377998 82170 378054 82226
rect 378122 82170 378178 82226
rect 378246 82170 378302 82226
rect 377874 82046 377930 82102
rect 377998 82046 378054 82102
rect 378122 82046 378178 82102
rect 378246 82046 378302 82102
rect 377874 81922 377930 81978
rect 377998 81922 378054 81978
rect 378122 81922 378178 81978
rect 378246 81922 378302 81978
rect 377874 64294 377930 64350
rect 377998 64294 378054 64350
rect 378122 64294 378178 64350
rect 378246 64294 378302 64350
rect 377874 64170 377930 64226
rect 377998 64170 378054 64226
rect 378122 64170 378178 64226
rect 378246 64170 378302 64226
rect 377874 64046 377930 64102
rect 377998 64046 378054 64102
rect 378122 64046 378178 64102
rect 378246 64046 378302 64102
rect 377874 63922 377930 63978
rect 377998 63922 378054 63978
rect 378122 63922 378178 63978
rect 378246 63922 378302 63978
rect 377874 46294 377930 46350
rect 377998 46294 378054 46350
rect 378122 46294 378178 46350
rect 378246 46294 378302 46350
rect 377874 46170 377930 46226
rect 377998 46170 378054 46226
rect 378122 46170 378178 46226
rect 378246 46170 378302 46226
rect 377874 46046 377930 46102
rect 377998 46046 378054 46102
rect 378122 46046 378178 46102
rect 378246 46046 378302 46102
rect 377874 45922 377930 45978
rect 377998 45922 378054 45978
rect 378122 45922 378178 45978
rect 378246 45922 378302 45978
rect 377874 28294 377930 28350
rect 377998 28294 378054 28350
rect 378122 28294 378178 28350
rect 378246 28294 378302 28350
rect 377874 28170 377930 28226
rect 377998 28170 378054 28226
rect 378122 28170 378178 28226
rect 378246 28170 378302 28226
rect 377874 28046 377930 28102
rect 377998 28046 378054 28102
rect 378122 28046 378178 28102
rect 378246 28046 378302 28102
rect 377874 27922 377930 27978
rect 377998 27922 378054 27978
rect 378122 27922 378178 27978
rect 378246 27922 378302 27978
rect 377874 10294 377930 10350
rect 377998 10294 378054 10350
rect 378122 10294 378178 10350
rect 378246 10294 378302 10350
rect 377874 10170 377930 10226
rect 377998 10170 378054 10226
rect 378122 10170 378178 10226
rect 378246 10170 378302 10226
rect 377874 10046 377930 10102
rect 377998 10046 378054 10102
rect 378122 10046 378178 10102
rect 378246 10046 378302 10102
rect 377874 9922 377930 9978
rect 377998 9922 378054 9978
rect 378122 9922 378178 9978
rect 378246 9922 378302 9978
rect 377874 -1176 377930 -1120
rect 377998 -1176 378054 -1120
rect 378122 -1176 378178 -1120
rect 378246 -1176 378302 -1120
rect 377874 -1300 377930 -1244
rect 377998 -1300 378054 -1244
rect 378122 -1300 378178 -1244
rect 378246 -1300 378302 -1244
rect 377874 -1424 377930 -1368
rect 377998 -1424 378054 -1368
rect 378122 -1424 378178 -1368
rect 378246 -1424 378302 -1368
rect 377874 -1548 377930 -1492
rect 377998 -1548 378054 -1492
rect 378122 -1548 378178 -1492
rect 378246 -1548 378302 -1492
rect 404874 130294 404930 130350
rect 404998 130294 405054 130350
rect 405122 130294 405178 130350
rect 405246 130294 405302 130350
rect 404874 130170 404930 130226
rect 404998 130170 405054 130226
rect 405122 130170 405178 130226
rect 405246 130170 405302 130226
rect 404874 130046 404930 130102
rect 404998 130046 405054 130102
rect 405122 130046 405178 130102
rect 405246 130046 405302 130102
rect 404874 129922 404930 129978
rect 404998 129922 405054 129978
rect 405122 129922 405178 129978
rect 405246 129922 405302 129978
rect 404874 112294 404930 112350
rect 404998 112294 405054 112350
rect 405122 112294 405178 112350
rect 405246 112294 405302 112350
rect 404874 112170 404930 112226
rect 404998 112170 405054 112226
rect 405122 112170 405178 112226
rect 405246 112170 405302 112226
rect 404874 112046 404930 112102
rect 404998 112046 405054 112102
rect 405122 112046 405178 112102
rect 405246 112046 405302 112102
rect 404874 111922 404930 111978
rect 404998 111922 405054 111978
rect 405122 111922 405178 111978
rect 405246 111922 405302 111978
rect 404874 94294 404930 94350
rect 404998 94294 405054 94350
rect 405122 94294 405178 94350
rect 405246 94294 405302 94350
rect 404874 94170 404930 94226
rect 404998 94170 405054 94226
rect 405122 94170 405178 94226
rect 405246 94170 405302 94226
rect 404874 94046 404930 94102
rect 404998 94046 405054 94102
rect 405122 94046 405178 94102
rect 405246 94046 405302 94102
rect 404874 93922 404930 93978
rect 404998 93922 405054 93978
rect 405122 93922 405178 93978
rect 405246 93922 405302 93978
rect 404874 76294 404930 76350
rect 404998 76294 405054 76350
rect 405122 76294 405178 76350
rect 405246 76294 405302 76350
rect 404874 76170 404930 76226
rect 404998 76170 405054 76226
rect 405122 76170 405178 76226
rect 405246 76170 405302 76226
rect 404874 76046 404930 76102
rect 404998 76046 405054 76102
rect 405122 76046 405178 76102
rect 405246 76046 405302 76102
rect 404874 75922 404930 75978
rect 404998 75922 405054 75978
rect 405122 75922 405178 75978
rect 405246 75922 405302 75978
rect 404874 58294 404930 58350
rect 404998 58294 405054 58350
rect 405122 58294 405178 58350
rect 405246 58294 405302 58350
rect 404874 58170 404930 58226
rect 404998 58170 405054 58226
rect 405122 58170 405178 58226
rect 405246 58170 405302 58226
rect 404874 58046 404930 58102
rect 404998 58046 405054 58102
rect 405122 58046 405178 58102
rect 405246 58046 405302 58102
rect 404874 57922 404930 57978
rect 404998 57922 405054 57978
rect 405122 57922 405178 57978
rect 405246 57922 405302 57978
rect 404874 40294 404930 40350
rect 404998 40294 405054 40350
rect 405122 40294 405178 40350
rect 405246 40294 405302 40350
rect 404874 40170 404930 40226
rect 404998 40170 405054 40226
rect 405122 40170 405178 40226
rect 405246 40170 405302 40226
rect 404874 40046 404930 40102
rect 404998 40046 405054 40102
rect 405122 40046 405178 40102
rect 405246 40046 405302 40102
rect 404874 39922 404930 39978
rect 404998 39922 405054 39978
rect 405122 39922 405178 39978
rect 405246 39922 405302 39978
rect 404874 22294 404930 22350
rect 404998 22294 405054 22350
rect 405122 22294 405178 22350
rect 405246 22294 405302 22350
rect 404874 22170 404930 22226
rect 404998 22170 405054 22226
rect 405122 22170 405178 22226
rect 405246 22170 405302 22226
rect 404874 22046 404930 22102
rect 404998 22046 405054 22102
rect 405122 22046 405178 22102
rect 405246 22046 405302 22102
rect 404874 21922 404930 21978
rect 404998 21922 405054 21978
rect 405122 21922 405178 21978
rect 405246 21922 405302 21978
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 408594 388294 408650 388350
rect 408718 388294 408774 388350
rect 408842 388294 408898 388350
rect 408966 388294 409022 388350
rect 408594 388170 408650 388226
rect 408718 388170 408774 388226
rect 408842 388170 408898 388226
rect 408966 388170 409022 388226
rect 408594 388046 408650 388102
rect 408718 388046 408774 388102
rect 408842 388046 408898 388102
rect 408966 388046 409022 388102
rect 408594 387922 408650 387978
rect 408718 387922 408774 387978
rect 408842 387922 408898 387978
rect 408966 387922 409022 387978
rect 408594 370294 408650 370350
rect 408718 370294 408774 370350
rect 408842 370294 408898 370350
rect 408966 370294 409022 370350
rect 408594 370170 408650 370226
rect 408718 370170 408774 370226
rect 408842 370170 408898 370226
rect 408966 370170 409022 370226
rect 408594 370046 408650 370102
rect 408718 370046 408774 370102
rect 408842 370046 408898 370102
rect 408966 370046 409022 370102
rect 408594 369922 408650 369978
rect 408718 369922 408774 369978
rect 408842 369922 408898 369978
rect 408966 369922 409022 369978
rect 408594 352294 408650 352350
rect 408718 352294 408774 352350
rect 408842 352294 408898 352350
rect 408966 352294 409022 352350
rect 408594 352170 408650 352226
rect 408718 352170 408774 352226
rect 408842 352170 408898 352226
rect 408966 352170 409022 352226
rect 408594 352046 408650 352102
rect 408718 352046 408774 352102
rect 408842 352046 408898 352102
rect 408966 352046 409022 352102
rect 408594 351922 408650 351978
rect 408718 351922 408774 351978
rect 408842 351922 408898 351978
rect 408966 351922 409022 351978
rect 408594 334294 408650 334350
rect 408718 334294 408774 334350
rect 408842 334294 408898 334350
rect 408966 334294 409022 334350
rect 408594 334170 408650 334226
rect 408718 334170 408774 334226
rect 408842 334170 408898 334226
rect 408966 334170 409022 334226
rect 408594 334046 408650 334102
rect 408718 334046 408774 334102
rect 408842 334046 408898 334102
rect 408966 334046 409022 334102
rect 408594 333922 408650 333978
rect 408718 333922 408774 333978
rect 408842 333922 408898 333978
rect 408966 333922 409022 333978
rect 408594 316294 408650 316350
rect 408718 316294 408774 316350
rect 408842 316294 408898 316350
rect 408966 316294 409022 316350
rect 408594 316170 408650 316226
rect 408718 316170 408774 316226
rect 408842 316170 408898 316226
rect 408966 316170 409022 316226
rect 408594 316046 408650 316102
rect 408718 316046 408774 316102
rect 408842 316046 408898 316102
rect 408966 316046 409022 316102
rect 408594 315922 408650 315978
rect 408718 315922 408774 315978
rect 408842 315922 408898 315978
rect 408966 315922 409022 315978
rect 408594 298294 408650 298350
rect 408718 298294 408774 298350
rect 408842 298294 408898 298350
rect 408966 298294 409022 298350
rect 408594 298170 408650 298226
rect 408718 298170 408774 298226
rect 408842 298170 408898 298226
rect 408966 298170 409022 298226
rect 408594 298046 408650 298102
rect 408718 298046 408774 298102
rect 408842 298046 408898 298102
rect 408966 298046 409022 298102
rect 408594 297922 408650 297978
rect 408718 297922 408774 297978
rect 408842 297922 408898 297978
rect 408966 297922 409022 297978
rect 408594 280294 408650 280350
rect 408718 280294 408774 280350
rect 408842 280294 408898 280350
rect 408966 280294 409022 280350
rect 408594 280170 408650 280226
rect 408718 280170 408774 280226
rect 408842 280170 408898 280226
rect 408966 280170 409022 280226
rect 408594 280046 408650 280102
rect 408718 280046 408774 280102
rect 408842 280046 408898 280102
rect 408966 280046 409022 280102
rect 408594 279922 408650 279978
rect 408718 279922 408774 279978
rect 408842 279922 408898 279978
rect 408966 279922 409022 279978
rect 408594 262294 408650 262350
rect 408718 262294 408774 262350
rect 408842 262294 408898 262350
rect 408966 262294 409022 262350
rect 408594 262170 408650 262226
rect 408718 262170 408774 262226
rect 408842 262170 408898 262226
rect 408966 262170 409022 262226
rect 408594 262046 408650 262102
rect 408718 262046 408774 262102
rect 408842 262046 408898 262102
rect 408966 262046 409022 262102
rect 408594 261922 408650 261978
rect 408718 261922 408774 261978
rect 408842 261922 408898 261978
rect 408966 261922 409022 261978
rect 435594 400294 435650 400350
rect 435718 400294 435774 400350
rect 435842 400294 435898 400350
rect 435966 400294 436022 400350
rect 435594 400170 435650 400226
rect 435718 400170 435774 400226
rect 435842 400170 435898 400226
rect 435966 400170 436022 400226
rect 435594 400046 435650 400102
rect 435718 400046 435774 400102
rect 435842 400046 435898 400102
rect 435966 400046 436022 400102
rect 435594 399922 435650 399978
rect 435718 399922 435774 399978
rect 435842 399922 435898 399978
rect 435966 399922 436022 399978
rect 435594 382294 435650 382350
rect 435718 382294 435774 382350
rect 435842 382294 435898 382350
rect 435966 382294 436022 382350
rect 435594 382170 435650 382226
rect 435718 382170 435774 382226
rect 435842 382170 435898 382226
rect 435966 382170 436022 382226
rect 435594 382046 435650 382102
rect 435718 382046 435774 382102
rect 435842 382046 435898 382102
rect 435966 382046 436022 382102
rect 435594 381922 435650 381978
rect 435718 381922 435774 381978
rect 435842 381922 435898 381978
rect 435966 381922 436022 381978
rect 435594 364294 435650 364350
rect 435718 364294 435774 364350
rect 435842 364294 435898 364350
rect 435966 364294 436022 364350
rect 435594 364170 435650 364226
rect 435718 364170 435774 364226
rect 435842 364170 435898 364226
rect 435966 364170 436022 364226
rect 435594 364046 435650 364102
rect 435718 364046 435774 364102
rect 435842 364046 435898 364102
rect 435966 364046 436022 364102
rect 435594 363922 435650 363978
rect 435718 363922 435774 363978
rect 435842 363922 435898 363978
rect 435966 363922 436022 363978
rect 435594 346294 435650 346350
rect 435718 346294 435774 346350
rect 435842 346294 435898 346350
rect 435966 346294 436022 346350
rect 435594 346170 435650 346226
rect 435718 346170 435774 346226
rect 435842 346170 435898 346226
rect 435966 346170 436022 346226
rect 435594 346046 435650 346102
rect 435718 346046 435774 346102
rect 435842 346046 435898 346102
rect 435966 346046 436022 346102
rect 435594 345922 435650 345978
rect 435718 345922 435774 345978
rect 435842 345922 435898 345978
rect 435966 345922 436022 345978
rect 435594 328294 435650 328350
rect 435718 328294 435774 328350
rect 435842 328294 435898 328350
rect 435966 328294 436022 328350
rect 435594 328170 435650 328226
rect 435718 328170 435774 328226
rect 435842 328170 435898 328226
rect 435966 328170 436022 328226
rect 435594 328046 435650 328102
rect 435718 328046 435774 328102
rect 435842 328046 435898 328102
rect 435966 328046 436022 328102
rect 435594 327922 435650 327978
rect 435718 327922 435774 327978
rect 435842 327922 435898 327978
rect 435966 327922 436022 327978
rect 435594 310294 435650 310350
rect 435718 310294 435774 310350
rect 435842 310294 435898 310350
rect 435966 310294 436022 310350
rect 435594 310170 435650 310226
rect 435718 310170 435774 310226
rect 435842 310170 435898 310226
rect 435966 310170 436022 310226
rect 435594 310046 435650 310102
rect 435718 310046 435774 310102
rect 435842 310046 435898 310102
rect 435966 310046 436022 310102
rect 435594 309922 435650 309978
rect 435718 309922 435774 309978
rect 435842 309922 435898 309978
rect 435966 309922 436022 309978
rect 435594 292294 435650 292350
rect 435718 292294 435774 292350
rect 435842 292294 435898 292350
rect 435966 292294 436022 292350
rect 435594 292170 435650 292226
rect 435718 292170 435774 292226
rect 435842 292170 435898 292226
rect 435966 292170 436022 292226
rect 435594 292046 435650 292102
rect 435718 292046 435774 292102
rect 435842 292046 435898 292102
rect 435966 292046 436022 292102
rect 435594 291922 435650 291978
rect 435718 291922 435774 291978
rect 435842 291922 435898 291978
rect 435966 291922 436022 291978
rect 435594 274294 435650 274350
rect 435718 274294 435774 274350
rect 435842 274294 435898 274350
rect 435966 274294 436022 274350
rect 435594 274170 435650 274226
rect 435718 274170 435774 274226
rect 435842 274170 435898 274226
rect 435966 274170 436022 274226
rect 435594 274046 435650 274102
rect 435718 274046 435774 274102
rect 435842 274046 435898 274102
rect 435966 274046 436022 274102
rect 435594 273922 435650 273978
rect 435718 273922 435774 273978
rect 435842 273922 435898 273978
rect 435966 273922 436022 273978
rect 408594 244294 408650 244350
rect 408718 244294 408774 244350
rect 408842 244294 408898 244350
rect 408966 244294 409022 244350
rect 408594 244170 408650 244226
rect 408718 244170 408774 244226
rect 408842 244170 408898 244226
rect 408966 244170 409022 244226
rect 408594 244046 408650 244102
rect 408718 244046 408774 244102
rect 408842 244046 408898 244102
rect 408966 244046 409022 244102
rect 408594 243922 408650 243978
rect 408718 243922 408774 243978
rect 408842 243922 408898 243978
rect 408966 243922 409022 243978
rect 408594 226294 408650 226350
rect 408718 226294 408774 226350
rect 408842 226294 408898 226350
rect 408966 226294 409022 226350
rect 408594 226170 408650 226226
rect 408718 226170 408774 226226
rect 408842 226170 408898 226226
rect 408966 226170 409022 226226
rect 408594 226046 408650 226102
rect 408718 226046 408774 226102
rect 408842 226046 408898 226102
rect 408966 226046 409022 226102
rect 408594 225922 408650 225978
rect 408718 225922 408774 225978
rect 408842 225922 408898 225978
rect 408966 225922 409022 225978
rect 408594 208294 408650 208350
rect 408718 208294 408774 208350
rect 408842 208294 408898 208350
rect 408966 208294 409022 208350
rect 408594 208170 408650 208226
rect 408718 208170 408774 208226
rect 408842 208170 408898 208226
rect 408966 208170 409022 208226
rect 408594 208046 408650 208102
rect 408718 208046 408774 208102
rect 408842 208046 408898 208102
rect 408966 208046 409022 208102
rect 408594 207922 408650 207978
rect 408718 207922 408774 207978
rect 408842 207922 408898 207978
rect 408966 207922 409022 207978
rect 408594 190294 408650 190350
rect 408718 190294 408774 190350
rect 408842 190294 408898 190350
rect 408966 190294 409022 190350
rect 408594 190170 408650 190226
rect 408718 190170 408774 190226
rect 408842 190170 408898 190226
rect 408966 190170 409022 190226
rect 408594 190046 408650 190102
rect 408718 190046 408774 190102
rect 408842 190046 408898 190102
rect 408966 190046 409022 190102
rect 408594 189922 408650 189978
rect 408718 189922 408774 189978
rect 408842 189922 408898 189978
rect 408966 189922 409022 189978
rect 408594 172294 408650 172350
rect 408718 172294 408774 172350
rect 408842 172294 408898 172350
rect 408966 172294 409022 172350
rect 408594 172170 408650 172226
rect 408718 172170 408774 172226
rect 408842 172170 408898 172226
rect 408966 172170 409022 172226
rect 408594 172046 408650 172102
rect 408718 172046 408774 172102
rect 408842 172046 408898 172102
rect 408966 172046 409022 172102
rect 408594 171922 408650 171978
rect 408718 171922 408774 171978
rect 408842 171922 408898 171978
rect 408966 171922 409022 171978
rect 408594 154294 408650 154350
rect 408718 154294 408774 154350
rect 408842 154294 408898 154350
rect 408966 154294 409022 154350
rect 408594 154170 408650 154226
rect 408718 154170 408774 154226
rect 408842 154170 408898 154226
rect 408966 154170 409022 154226
rect 408594 154046 408650 154102
rect 408718 154046 408774 154102
rect 408842 154046 408898 154102
rect 408966 154046 409022 154102
rect 408594 153922 408650 153978
rect 408718 153922 408774 153978
rect 408842 153922 408898 153978
rect 408966 153922 409022 153978
rect 418348 142622 418404 142678
rect 418348 141902 418404 141958
rect 414652 141002 414708 141058
rect 435594 256294 435650 256350
rect 435718 256294 435774 256350
rect 435842 256294 435898 256350
rect 435966 256294 436022 256350
rect 435594 256170 435650 256226
rect 435718 256170 435774 256226
rect 435842 256170 435898 256226
rect 435966 256170 436022 256226
rect 435594 256046 435650 256102
rect 435718 256046 435774 256102
rect 435842 256046 435898 256102
rect 435966 256046 436022 256102
rect 435594 255922 435650 255978
rect 435718 255922 435774 255978
rect 435842 255922 435898 255978
rect 435966 255922 436022 255978
rect 435594 238294 435650 238350
rect 435718 238294 435774 238350
rect 435842 238294 435898 238350
rect 435966 238294 436022 238350
rect 435594 238170 435650 238226
rect 435718 238170 435774 238226
rect 435842 238170 435898 238226
rect 435966 238170 436022 238226
rect 435594 238046 435650 238102
rect 435718 238046 435774 238102
rect 435842 238046 435898 238102
rect 435966 238046 436022 238102
rect 435594 237922 435650 237978
rect 435718 237922 435774 237978
rect 435842 237922 435898 237978
rect 435966 237922 436022 237978
rect 435594 220294 435650 220350
rect 435718 220294 435774 220350
rect 435842 220294 435898 220350
rect 435966 220294 436022 220350
rect 435594 220170 435650 220226
rect 435718 220170 435774 220226
rect 435842 220170 435898 220226
rect 435966 220170 436022 220226
rect 435594 220046 435650 220102
rect 435718 220046 435774 220102
rect 435842 220046 435898 220102
rect 435966 220046 436022 220102
rect 435594 219922 435650 219978
rect 435718 219922 435774 219978
rect 435842 219922 435898 219978
rect 435966 219922 436022 219978
rect 435594 202294 435650 202350
rect 435718 202294 435774 202350
rect 435842 202294 435898 202350
rect 435966 202294 436022 202350
rect 435594 202170 435650 202226
rect 435718 202170 435774 202226
rect 435842 202170 435898 202226
rect 435966 202170 436022 202226
rect 435594 202046 435650 202102
rect 435718 202046 435774 202102
rect 435842 202046 435898 202102
rect 435966 202046 436022 202102
rect 435594 201922 435650 201978
rect 435718 201922 435774 201978
rect 435842 201922 435898 201978
rect 435966 201922 436022 201978
rect 435594 184294 435650 184350
rect 435718 184294 435774 184350
rect 435842 184294 435898 184350
rect 435966 184294 436022 184350
rect 435594 184170 435650 184226
rect 435718 184170 435774 184226
rect 435842 184170 435898 184226
rect 435966 184170 436022 184226
rect 435594 184046 435650 184102
rect 435718 184046 435774 184102
rect 435842 184046 435898 184102
rect 435966 184046 436022 184102
rect 435594 183922 435650 183978
rect 435718 183922 435774 183978
rect 435842 183922 435898 183978
rect 435966 183922 436022 183978
rect 435594 166294 435650 166350
rect 435718 166294 435774 166350
rect 435842 166294 435898 166350
rect 435966 166294 436022 166350
rect 435594 166170 435650 166226
rect 435718 166170 435774 166226
rect 435842 166170 435898 166226
rect 435966 166170 436022 166226
rect 435594 166046 435650 166102
rect 435718 166046 435774 166102
rect 435842 166046 435898 166102
rect 435966 166046 436022 166102
rect 435594 165922 435650 165978
rect 435718 165922 435774 165978
rect 435842 165922 435898 165978
rect 435966 165922 436022 165978
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 408594 136294 408650 136350
rect 408718 136294 408774 136350
rect 408842 136294 408898 136350
rect 408966 136294 409022 136350
rect 408594 136170 408650 136226
rect 408718 136170 408774 136226
rect 408842 136170 408898 136226
rect 408966 136170 409022 136226
rect 408594 136046 408650 136102
rect 408718 136046 408774 136102
rect 408842 136046 408898 136102
rect 408966 136046 409022 136102
rect 408594 135922 408650 135978
rect 408718 135922 408774 135978
rect 408842 135922 408898 135978
rect 408966 135922 409022 135978
rect 408594 118294 408650 118350
rect 408718 118294 408774 118350
rect 408842 118294 408898 118350
rect 408966 118294 409022 118350
rect 408594 118170 408650 118226
rect 408718 118170 408774 118226
rect 408842 118170 408898 118226
rect 408966 118170 409022 118226
rect 408594 118046 408650 118102
rect 408718 118046 408774 118102
rect 408842 118046 408898 118102
rect 408966 118046 409022 118102
rect 408594 117922 408650 117978
rect 408718 117922 408774 117978
rect 408842 117922 408898 117978
rect 408966 117922 409022 117978
rect 408594 100294 408650 100350
rect 408718 100294 408774 100350
rect 408842 100294 408898 100350
rect 408966 100294 409022 100350
rect 408594 100170 408650 100226
rect 408718 100170 408774 100226
rect 408842 100170 408898 100226
rect 408966 100170 409022 100226
rect 408594 100046 408650 100102
rect 408718 100046 408774 100102
rect 408842 100046 408898 100102
rect 408966 100046 409022 100102
rect 408594 99922 408650 99978
rect 408718 99922 408774 99978
rect 408842 99922 408898 99978
rect 408966 99922 409022 99978
rect 408594 82294 408650 82350
rect 408718 82294 408774 82350
rect 408842 82294 408898 82350
rect 408966 82294 409022 82350
rect 408594 82170 408650 82226
rect 408718 82170 408774 82226
rect 408842 82170 408898 82226
rect 408966 82170 409022 82226
rect 408594 82046 408650 82102
rect 408718 82046 408774 82102
rect 408842 82046 408898 82102
rect 408966 82046 409022 82102
rect 408594 81922 408650 81978
rect 408718 81922 408774 81978
rect 408842 81922 408898 81978
rect 408966 81922 409022 81978
rect 408594 64294 408650 64350
rect 408718 64294 408774 64350
rect 408842 64294 408898 64350
rect 408966 64294 409022 64350
rect 408594 64170 408650 64226
rect 408718 64170 408774 64226
rect 408842 64170 408898 64226
rect 408966 64170 409022 64226
rect 408594 64046 408650 64102
rect 408718 64046 408774 64102
rect 408842 64046 408898 64102
rect 408966 64046 409022 64102
rect 408594 63922 408650 63978
rect 408718 63922 408774 63978
rect 408842 63922 408898 63978
rect 408966 63922 409022 63978
rect 408594 46294 408650 46350
rect 408718 46294 408774 46350
rect 408842 46294 408898 46350
rect 408966 46294 409022 46350
rect 408594 46170 408650 46226
rect 408718 46170 408774 46226
rect 408842 46170 408898 46226
rect 408966 46170 409022 46226
rect 408594 46046 408650 46102
rect 408718 46046 408774 46102
rect 408842 46046 408898 46102
rect 408966 46046 409022 46102
rect 408594 45922 408650 45978
rect 408718 45922 408774 45978
rect 408842 45922 408898 45978
rect 408966 45922 409022 45978
rect 408594 28294 408650 28350
rect 408718 28294 408774 28350
rect 408842 28294 408898 28350
rect 408966 28294 409022 28350
rect 408594 28170 408650 28226
rect 408718 28170 408774 28226
rect 408842 28170 408898 28226
rect 408966 28170 409022 28226
rect 408594 28046 408650 28102
rect 408718 28046 408774 28102
rect 408842 28046 408898 28102
rect 408966 28046 409022 28102
rect 408594 27922 408650 27978
rect 408718 27922 408774 27978
rect 408842 27922 408898 27978
rect 408966 27922 409022 27978
rect 408594 10294 408650 10350
rect 408718 10294 408774 10350
rect 408842 10294 408898 10350
rect 408966 10294 409022 10350
rect 408594 10170 408650 10226
rect 408718 10170 408774 10226
rect 408842 10170 408898 10226
rect 408966 10170 409022 10226
rect 408594 10046 408650 10102
rect 408718 10046 408774 10102
rect 408842 10046 408898 10102
rect 408966 10046 409022 10102
rect 408594 9922 408650 9978
rect 408718 9922 408774 9978
rect 408842 9922 408898 9978
rect 408966 9922 409022 9978
rect 408594 -1176 408650 -1120
rect 408718 -1176 408774 -1120
rect 408842 -1176 408898 -1120
rect 408966 -1176 409022 -1120
rect 408594 -1300 408650 -1244
rect 408718 -1300 408774 -1244
rect 408842 -1300 408898 -1244
rect 408966 -1300 409022 -1244
rect 408594 -1424 408650 -1368
rect 408718 -1424 408774 -1368
rect 408842 -1424 408898 -1368
rect 408966 -1424 409022 -1368
rect 408594 -1548 408650 -1492
rect 408718 -1548 408774 -1492
rect 408842 -1548 408898 -1492
rect 408966 -1548 409022 -1492
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 439314 388294 439370 388350
rect 439438 388294 439494 388350
rect 439562 388294 439618 388350
rect 439686 388294 439742 388350
rect 439314 388170 439370 388226
rect 439438 388170 439494 388226
rect 439562 388170 439618 388226
rect 439686 388170 439742 388226
rect 439314 388046 439370 388102
rect 439438 388046 439494 388102
rect 439562 388046 439618 388102
rect 439686 388046 439742 388102
rect 439314 387922 439370 387978
rect 439438 387922 439494 387978
rect 439562 387922 439618 387978
rect 439686 387922 439742 387978
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 470034 568294 470090 568350
rect 470158 568294 470214 568350
rect 470282 568294 470338 568350
rect 470406 568294 470462 568350
rect 470034 568170 470090 568226
rect 470158 568170 470214 568226
rect 470282 568170 470338 568226
rect 470406 568170 470462 568226
rect 470034 568046 470090 568102
rect 470158 568046 470214 568102
rect 470282 568046 470338 568102
rect 470406 568046 470462 568102
rect 470034 567922 470090 567978
rect 470158 567922 470214 567978
rect 470282 567922 470338 567978
rect 470406 567922 470462 567978
rect 470034 550294 470090 550350
rect 470158 550294 470214 550350
rect 470282 550294 470338 550350
rect 470406 550294 470462 550350
rect 470034 550170 470090 550226
rect 470158 550170 470214 550226
rect 470282 550170 470338 550226
rect 470406 550170 470462 550226
rect 470034 550046 470090 550102
rect 470158 550046 470214 550102
rect 470282 550046 470338 550102
rect 470406 550046 470462 550102
rect 470034 549922 470090 549978
rect 470158 549922 470214 549978
rect 470282 549922 470338 549978
rect 470406 549922 470462 549978
rect 466314 544294 466370 544350
rect 466438 544294 466494 544350
rect 466562 544294 466618 544350
rect 466686 544294 466742 544350
rect 466314 544170 466370 544226
rect 466438 544170 466494 544226
rect 466562 544170 466618 544226
rect 466686 544170 466742 544226
rect 466314 544046 466370 544102
rect 466438 544046 466494 544102
rect 466562 544046 466618 544102
rect 466686 544046 466742 544102
rect 466314 543922 466370 543978
rect 466438 543922 466494 543978
rect 466562 543922 466618 543978
rect 466686 543922 466742 543978
rect 466314 526294 466370 526350
rect 466438 526294 466494 526350
rect 466562 526294 466618 526350
rect 466686 526294 466742 526350
rect 466314 526170 466370 526226
rect 466438 526170 466494 526226
rect 466562 526170 466618 526226
rect 466686 526170 466742 526226
rect 466314 526046 466370 526102
rect 466438 526046 466494 526102
rect 466562 526046 466618 526102
rect 466686 526046 466742 526102
rect 466314 525922 466370 525978
rect 466438 525922 466494 525978
rect 466562 525922 466618 525978
rect 466686 525922 466742 525978
rect 466314 508294 466370 508350
rect 466438 508294 466494 508350
rect 466562 508294 466618 508350
rect 466686 508294 466742 508350
rect 466314 508170 466370 508226
rect 466438 508170 466494 508226
rect 466562 508170 466618 508226
rect 466686 508170 466742 508226
rect 466314 508046 466370 508102
rect 466438 508046 466494 508102
rect 466562 508046 466618 508102
rect 466686 508046 466742 508102
rect 466314 507922 466370 507978
rect 466438 507922 466494 507978
rect 466562 507922 466618 507978
rect 466686 507922 466742 507978
rect 466314 490294 466370 490350
rect 466438 490294 466494 490350
rect 466562 490294 466618 490350
rect 466686 490294 466742 490350
rect 466314 490170 466370 490226
rect 466438 490170 466494 490226
rect 466562 490170 466618 490226
rect 466686 490170 466742 490226
rect 466314 490046 466370 490102
rect 466438 490046 466494 490102
rect 466562 490046 466618 490102
rect 466686 490046 466742 490102
rect 466314 489922 466370 489978
rect 466438 489922 466494 489978
rect 466562 489922 466618 489978
rect 466686 489922 466742 489978
rect 470034 532294 470090 532350
rect 470158 532294 470214 532350
rect 470282 532294 470338 532350
rect 470406 532294 470462 532350
rect 470034 532170 470090 532226
rect 470158 532170 470214 532226
rect 470282 532170 470338 532226
rect 470406 532170 470462 532226
rect 470034 532046 470090 532102
rect 470158 532046 470214 532102
rect 470282 532046 470338 532102
rect 470406 532046 470462 532102
rect 470034 531922 470090 531978
rect 470158 531922 470214 531978
rect 470282 531922 470338 531978
rect 470406 531922 470462 531978
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 497034 562294 497090 562350
rect 497158 562294 497214 562350
rect 497282 562294 497338 562350
rect 497406 562294 497462 562350
rect 497034 562170 497090 562226
rect 497158 562170 497214 562226
rect 497282 562170 497338 562226
rect 497406 562170 497462 562226
rect 497034 562046 497090 562102
rect 497158 562046 497214 562102
rect 497282 562046 497338 562102
rect 497406 562046 497462 562102
rect 497034 561922 497090 561978
rect 497158 561922 497214 561978
rect 497282 561922 497338 561978
rect 497406 561922 497462 561978
rect 497034 544294 497090 544350
rect 497158 544294 497214 544350
rect 497282 544294 497338 544350
rect 497406 544294 497462 544350
rect 497034 544170 497090 544226
rect 497158 544170 497214 544226
rect 497282 544170 497338 544226
rect 497406 544170 497462 544226
rect 497034 544046 497090 544102
rect 497158 544046 497214 544102
rect 497282 544046 497338 544102
rect 497406 544046 497462 544102
rect 497034 543922 497090 543978
rect 497158 543922 497214 543978
rect 497282 543922 497338 543978
rect 497406 543922 497462 543978
rect 474518 526294 474574 526350
rect 474642 526294 474698 526350
rect 497034 526376 497090 526432
rect 497158 526376 497214 526432
rect 497282 526376 497338 526432
rect 497406 526376 497462 526432
rect 497034 526252 497090 526308
rect 497158 526252 497214 526308
rect 497282 526252 497338 526308
rect 497406 526252 497462 526308
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 500754 568294 500810 568350
rect 500878 568294 500934 568350
rect 501002 568294 501058 568350
rect 501126 568294 501182 568350
rect 500754 568170 500810 568226
rect 500878 568170 500934 568226
rect 501002 568170 501058 568226
rect 501126 568170 501182 568226
rect 500754 568046 500810 568102
rect 500878 568046 500934 568102
rect 501002 568046 501058 568102
rect 501126 568046 501182 568102
rect 500754 567922 500810 567978
rect 500878 567922 500934 567978
rect 501002 567922 501058 567978
rect 501126 567922 501182 567978
rect 500754 550294 500810 550350
rect 500878 550294 500934 550350
rect 501002 550294 501058 550350
rect 501126 550294 501182 550350
rect 500754 550170 500810 550226
rect 500878 550170 500934 550226
rect 501002 550170 501058 550226
rect 501126 550170 501182 550226
rect 500754 550046 500810 550102
rect 500878 550046 500934 550102
rect 501002 550046 501058 550102
rect 501126 550046 501182 550102
rect 500754 549922 500810 549978
rect 500878 549922 500934 549978
rect 501002 549922 501058 549978
rect 501126 549922 501182 549978
rect 500754 532294 500810 532350
rect 500878 532294 500934 532350
rect 501002 532294 501058 532350
rect 501126 532294 501182 532350
rect 500754 532170 500810 532226
rect 500878 532170 500934 532226
rect 501002 532170 501058 532226
rect 501126 532170 501182 532226
rect 500754 532046 500810 532102
rect 500878 532046 500934 532102
rect 501002 532046 501058 532102
rect 501126 532046 501182 532102
rect 500754 531922 500810 531978
rect 500878 531922 500934 531978
rect 501002 531922 501058 531978
rect 501126 531922 501182 531978
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 527754 562294 527810 562350
rect 527878 562294 527934 562350
rect 528002 562294 528058 562350
rect 528126 562294 528182 562350
rect 527754 562170 527810 562226
rect 527878 562170 527934 562226
rect 528002 562170 528058 562226
rect 528126 562170 528182 562226
rect 527754 562046 527810 562102
rect 527878 562046 527934 562102
rect 528002 562046 528058 562102
rect 528126 562046 528182 562102
rect 527754 561922 527810 561978
rect 527878 561922 527934 561978
rect 528002 561922 528058 561978
rect 528126 561922 528182 561978
rect 527754 544294 527810 544350
rect 527878 544294 527934 544350
rect 528002 544294 528058 544350
rect 528126 544294 528182 544350
rect 527754 544170 527810 544226
rect 527878 544170 527934 544226
rect 528002 544170 528058 544226
rect 528126 544170 528182 544226
rect 527754 544046 527810 544102
rect 527878 544046 527934 544102
rect 528002 544046 528058 544102
rect 528126 544046 528182 544102
rect 527754 543922 527810 543978
rect 527878 543922 527934 543978
rect 528002 543922 528058 543978
rect 528126 543922 528182 543978
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 531474 568294 531530 568350
rect 531598 568294 531654 568350
rect 531722 568294 531778 568350
rect 531846 568294 531902 568350
rect 531474 568170 531530 568226
rect 531598 568170 531654 568226
rect 531722 568170 531778 568226
rect 531846 568170 531902 568226
rect 531474 568046 531530 568102
rect 531598 568046 531654 568102
rect 531722 568046 531778 568102
rect 531846 568046 531902 568102
rect 531474 567922 531530 567978
rect 531598 567922 531654 567978
rect 531722 567922 531778 567978
rect 531846 567922 531902 567978
rect 531474 550294 531530 550350
rect 531598 550294 531654 550350
rect 531722 550294 531778 550350
rect 531846 550294 531902 550350
rect 531474 550170 531530 550226
rect 531598 550170 531654 550226
rect 531722 550170 531778 550226
rect 531846 550170 531902 550226
rect 531474 550046 531530 550102
rect 531598 550046 531654 550102
rect 531722 550046 531778 550102
rect 531846 550046 531902 550102
rect 531474 549922 531530 549978
rect 531598 549922 531654 549978
rect 531722 549922 531778 549978
rect 531846 549922 531902 549978
rect 505238 526294 505294 526350
rect 505362 526294 505418 526350
rect 474518 526170 474574 526226
rect 474642 526170 474698 526226
rect 474518 526046 474574 526102
rect 474642 526046 474698 526102
rect 474518 525922 474574 525978
rect 474642 525922 474698 525978
rect 527754 526376 527810 526432
rect 527878 526376 527934 526432
rect 528002 526376 528058 526432
rect 528126 526376 528182 526432
rect 527754 526252 527810 526308
rect 527878 526252 527934 526308
rect 528002 526252 528058 526308
rect 528126 526252 528182 526308
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 556220 546362 556276 546418
rect 556108 546182 556164 546238
rect 531474 532294 531530 532350
rect 531598 532294 531654 532350
rect 531722 532294 531778 532350
rect 531846 532294 531902 532350
rect 531474 532170 531530 532226
rect 531598 532170 531654 532226
rect 531722 532170 531778 532226
rect 531846 532170 531902 532226
rect 531474 532046 531530 532102
rect 531598 532046 531654 532102
rect 531722 532046 531778 532102
rect 531846 532046 531902 532102
rect 531474 531922 531530 531978
rect 531598 531922 531654 531978
rect 531722 531922 531778 531978
rect 531846 531922 531902 531978
rect 535958 526294 536014 526350
rect 536082 526294 536138 526350
rect 505238 526170 505294 526226
rect 505362 526170 505418 526226
rect 505238 526046 505294 526102
rect 505362 526046 505418 526102
rect 505238 525922 505294 525978
rect 505362 525922 505418 525978
rect 535958 526170 536014 526226
rect 536082 526170 536138 526226
rect 535958 526046 536014 526102
rect 536082 526046 536138 526102
rect 535958 525922 536014 525978
rect 536082 525922 536138 525978
rect 470034 514294 470090 514350
rect 470158 514294 470214 514350
rect 470282 514294 470338 514350
rect 470406 514294 470462 514350
rect 470034 514170 470090 514226
rect 470158 514170 470214 514226
rect 470282 514170 470338 514226
rect 470406 514170 470462 514226
rect 466314 472294 466370 472350
rect 466438 472294 466494 472350
rect 466562 472294 466618 472350
rect 466686 472294 466742 472350
rect 466314 472170 466370 472226
rect 466438 472170 466494 472226
rect 466562 472170 466618 472226
rect 466686 472170 466742 472226
rect 466314 472046 466370 472102
rect 466438 472046 466494 472102
rect 466562 472046 466618 472102
rect 466686 472046 466742 472102
rect 466314 471922 466370 471978
rect 466438 471922 466494 471978
rect 466562 471922 466618 471978
rect 466686 471922 466742 471978
rect 466314 454294 466370 454350
rect 466438 454294 466494 454350
rect 466562 454294 466618 454350
rect 466686 454294 466742 454350
rect 466314 454170 466370 454226
rect 466438 454170 466494 454226
rect 466562 454170 466618 454226
rect 466686 454170 466742 454226
rect 466314 454046 466370 454102
rect 466438 454046 466494 454102
rect 466562 454046 466618 454102
rect 466686 454046 466742 454102
rect 466314 453922 466370 453978
rect 466438 453922 466494 453978
rect 466562 453922 466618 453978
rect 466686 453922 466742 453978
rect 466314 436294 466370 436350
rect 466438 436294 466494 436350
rect 466562 436294 466618 436350
rect 466686 436294 466742 436350
rect 466314 436170 466370 436226
rect 466438 436170 466494 436226
rect 466562 436170 466618 436226
rect 466686 436170 466742 436226
rect 466314 436046 466370 436102
rect 466438 436046 466494 436102
rect 466562 436046 466618 436102
rect 466686 436046 466742 436102
rect 466314 435922 466370 435978
rect 466438 435922 466494 435978
rect 466562 435922 466618 435978
rect 466686 435922 466742 435978
rect 439314 370294 439370 370350
rect 439438 370294 439494 370350
rect 439562 370294 439618 370350
rect 439686 370294 439742 370350
rect 439314 370170 439370 370226
rect 439438 370170 439494 370226
rect 439562 370170 439618 370226
rect 439686 370170 439742 370226
rect 439314 370046 439370 370102
rect 439438 370046 439494 370102
rect 439562 370046 439618 370102
rect 439686 370046 439742 370102
rect 439314 369922 439370 369978
rect 439438 369922 439494 369978
rect 439562 369922 439618 369978
rect 439686 369922 439742 369978
rect 451164 371402 451220 371458
rect 451052 364742 451108 364798
rect 439314 352294 439370 352350
rect 439438 352294 439494 352350
rect 439562 352294 439618 352350
rect 439686 352294 439742 352350
rect 439314 352170 439370 352226
rect 439438 352170 439494 352226
rect 439562 352170 439618 352226
rect 439686 352170 439742 352226
rect 439314 352046 439370 352102
rect 439438 352046 439494 352102
rect 439562 352046 439618 352102
rect 439686 352046 439742 352102
rect 439314 351922 439370 351978
rect 439438 351922 439494 351978
rect 439562 351922 439618 351978
rect 439686 351922 439742 351978
rect 449484 354482 449540 354538
rect 449372 343502 449428 343558
rect 439314 334294 439370 334350
rect 439438 334294 439494 334350
rect 439562 334294 439618 334350
rect 439686 334294 439742 334350
rect 439314 334170 439370 334226
rect 439438 334170 439494 334226
rect 439562 334170 439618 334226
rect 439686 334170 439742 334226
rect 439314 334046 439370 334102
rect 439438 334046 439494 334102
rect 439562 334046 439618 334102
rect 439686 334046 439742 334102
rect 439314 333922 439370 333978
rect 439438 333922 439494 333978
rect 439562 333922 439618 333978
rect 439686 333922 439742 333978
rect 439314 316294 439370 316350
rect 439438 316294 439494 316350
rect 439562 316294 439618 316350
rect 439686 316294 439742 316350
rect 439314 316170 439370 316226
rect 439438 316170 439494 316226
rect 439562 316170 439618 316226
rect 439686 316170 439742 316226
rect 439314 316046 439370 316102
rect 439438 316046 439494 316102
rect 439562 316046 439618 316102
rect 439686 316046 439742 316102
rect 439314 315922 439370 315978
rect 439438 315922 439494 315978
rect 439562 315922 439618 315978
rect 439686 315922 439742 315978
rect 439314 298294 439370 298350
rect 439438 298294 439494 298350
rect 439562 298294 439618 298350
rect 439686 298294 439742 298350
rect 439314 298170 439370 298226
rect 439438 298170 439494 298226
rect 439562 298170 439618 298226
rect 439686 298170 439742 298226
rect 439314 298046 439370 298102
rect 439438 298046 439494 298102
rect 439562 298046 439618 298102
rect 439686 298046 439742 298102
rect 439314 297922 439370 297978
rect 439438 297922 439494 297978
rect 439562 297922 439618 297978
rect 439686 297922 439742 297978
rect 439314 280294 439370 280350
rect 439438 280294 439494 280350
rect 439562 280294 439618 280350
rect 439686 280294 439742 280350
rect 439314 280170 439370 280226
rect 439438 280170 439494 280226
rect 439562 280170 439618 280226
rect 439686 280170 439742 280226
rect 439314 280046 439370 280102
rect 439438 280046 439494 280102
rect 439562 280046 439618 280102
rect 439686 280046 439742 280102
rect 439314 279922 439370 279978
rect 439438 279922 439494 279978
rect 439562 279922 439618 279978
rect 439686 279922 439742 279978
rect 439314 262294 439370 262350
rect 439438 262294 439494 262350
rect 439562 262294 439618 262350
rect 439686 262294 439742 262350
rect 439314 262170 439370 262226
rect 439438 262170 439494 262226
rect 439562 262170 439618 262226
rect 439686 262170 439742 262226
rect 439314 262046 439370 262102
rect 439438 262046 439494 262102
rect 439562 262046 439618 262102
rect 439686 262046 439742 262102
rect 439314 261922 439370 261978
rect 439438 261922 439494 261978
rect 439562 261922 439618 261978
rect 439686 261922 439742 261978
rect 447468 341882 447524 341938
rect 439314 244294 439370 244350
rect 439438 244294 439494 244350
rect 439562 244294 439618 244350
rect 439686 244294 439742 244350
rect 439314 244170 439370 244226
rect 439438 244170 439494 244226
rect 439562 244170 439618 244226
rect 439686 244170 439742 244226
rect 439314 244046 439370 244102
rect 439438 244046 439494 244102
rect 439562 244046 439618 244102
rect 439686 244046 439742 244102
rect 439314 243922 439370 243978
rect 439438 243922 439494 243978
rect 439562 243922 439618 243978
rect 439686 243922 439742 243978
rect 439314 226294 439370 226350
rect 439438 226294 439494 226350
rect 439562 226294 439618 226350
rect 439686 226294 439742 226350
rect 439314 226170 439370 226226
rect 439438 226170 439494 226226
rect 439562 226170 439618 226226
rect 439686 226170 439742 226226
rect 439314 226046 439370 226102
rect 439438 226046 439494 226102
rect 439562 226046 439618 226102
rect 439686 226046 439742 226102
rect 439314 225922 439370 225978
rect 439438 225922 439494 225978
rect 439562 225922 439618 225978
rect 439686 225922 439742 225978
rect 439314 208294 439370 208350
rect 439438 208294 439494 208350
rect 439562 208294 439618 208350
rect 439686 208294 439742 208350
rect 439314 208170 439370 208226
rect 439438 208170 439494 208226
rect 439562 208170 439618 208226
rect 439686 208170 439742 208226
rect 439314 208046 439370 208102
rect 439438 208046 439494 208102
rect 439562 208046 439618 208102
rect 439686 208046 439742 208102
rect 439314 207922 439370 207978
rect 439438 207922 439494 207978
rect 439562 207922 439618 207978
rect 439686 207922 439742 207978
rect 439314 190294 439370 190350
rect 439438 190294 439494 190350
rect 439562 190294 439618 190350
rect 439686 190294 439742 190350
rect 439314 190170 439370 190226
rect 439438 190170 439494 190226
rect 439562 190170 439618 190226
rect 439686 190170 439742 190226
rect 439314 190046 439370 190102
rect 439438 190046 439494 190102
rect 439562 190046 439618 190102
rect 439686 190046 439742 190102
rect 439314 189922 439370 189978
rect 439438 189922 439494 189978
rect 439562 189922 439618 189978
rect 439686 189922 439742 189978
rect 439314 172294 439370 172350
rect 439438 172294 439494 172350
rect 439562 172294 439618 172350
rect 439686 172294 439742 172350
rect 439314 172170 439370 172226
rect 439438 172170 439494 172226
rect 439562 172170 439618 172226
rect 439686 172170 439742 172226
rect 439314 172046 439370 172102
rect 439438 172046 439494 172102
rect 439562 172046 439618 172102
rect 439686 172046 439742 172102
rect 439314 171922 439370 171978
rect 439438 171922 439494 171978
rect 439562 171922 439618 171978
rect 439686 171922 439742 171978
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 444668 142442 444724 142498
rect 446612 244294 446668 244350
rect 446736 244294 446792 244350
rect 446860 244294 446916 244350
rect 446984 244294 447040 244350
rect 446612 244170 446668 244226
rect 446736 244170 446792 244226
rect 446860 244170 446916 244226
rect 446984 244170 447040 244226
rect 446612 244046 446668 244102
rect 446736 244046 446792 244102
rect 446860 244046 446916 244102
rect 446984 244046 447040 244102
rect 446612 243922 446668 243978
rect 446736 243922 446792 243978
rect 446860 243922 446916 243978
rect 446984 243922 447040 243978
rect 445812 238294 445868 238350
rect 445936 238294 445992 238350
rect 446060 238294 446116 238350
rect 446184 238294 446240 238350
rect 445812 238170 445868 238226
rect 445936 238170 445992 238226
rect 446060 238170 446116 238226
rect 446184 238170 446240 238226
rect 445812 238046 445868 238102
rect 445936 238046 445992 238102
rect 446060 238046 446116 238102
rect 446184 238046 446240 238102
rect 445812 237922 445868 237978
rect 445936 237922 445992 237978
rect 446060 237922 446116 237978
rect 446184 237922 446240 237978
rect 446612 226294 446668 226350
rect 446736 226294 446792 226350
rect 446860 226294 446916 226350
rect 446984 226294 447040 226350
rect 446612 226170 446668 226226
rect 446736 226170 446792 226226
rect 446860 226170 446916 226226
rect 446984 226170 447040 226226
rect 446612 226046 446668 226102
rect 446736 226046 446792 226102
rect 446860 226046 446916 226102
rect 446984 226046 447040 226102
rect 446612 225922 446668 225978
rect 446736 225922 446792 225978
rect 446860 225922 446916 225978
rect 446984 225922 447040 225978
rect 445812 220294 445868 220350
rect 445936 220294 445992 220350
rect 446060 220294 446116 220350
rect 446184 220294 446240 220350
rect 445812 220170 445868 220226
rect 445936 220170 445992 220226
rect 446060 220170 446116 220226
rect 446184 220170 446240 220226
rect 445812 220046 445868 220102
rect 445936 220046 445992 220102
rect 446060 220046 446116 220102
rect 446184 220046 446240 220102
rect 445812 219922 445868 219978
rect 445936 219922 445992 219978
rect 446060 219922 446116 219978
rect 446184 219922 446240 219978
rect 446612 208294 446668 208350
rect 446736 208294 446792 208350
rect 446860 208294 446916 208350
rect 446984 208294 447040 208350
rect 446612 208170 446668 208226
rect 446736 208170 446792 208226
rect 446860 208170 446916 208226
rect 446984 208170 447040 208226
rect 446612 208046 446668 208102
rect 446736 208046 446792 208102
rect 446860 208046 446916 208102
rect 446984 208046 447040 208102
rect 446612 207922 446668 207978
rect 446736 207922 446792 207978
rect 446860 207922 446916 207978
rect 446984 207922 447040 207978
rect 445812 202294 445868 202350
rect 445936 202294 445992 202350
rect 446060 202294 446116 202350
rect 446184 202294 446240 202350
rect 445812 202170 445868 202226
rect 445936 202170 445992 202226
rect 446060 202170 446116 202226
rect 446184 202170 446240 202226
rect 445812 202046 445868 202102
rect 445936 202046 445992 202102
rect 446060 202046 446116 202102
rect 446184 202046 446240 202102
rect 445812 201922 445868 201978
rect 445936 201922 445992 201978
rect 446060 201922 446116 201978
rect 446184 201922 446240 201978
rect 446612 190294 446668 190350
rect 446736 190294 446792 190350
rect 446860 190294 446916 190350
rect 446984 190294 447040 190350
rect 446612 190170 446668 190226
rect 446736 190170 446792 190226
rect 446860 190170 446916 190226
rect 446984 190170 447040 190226
rect 446612 190046 446668 190102
rect 446736 190046 446792 190102
rect 446860 190046 446916 190102
rect 446984 190046 447040 190102
rect 446612 189922 446668 189978
rect 446736 189922 446792 189978
rect 446860 189922 446916 189978
rect 446984 189922 447040 189978
rect 445812 184294 445868 184350
rect 445936 184294 445992 184350
rect 446060 184294 446116 184350
rect 446184 184294 446240 184350
rect 445812 184170 445868 184226
rect 445936 184170 445992 184226
rect 446060 184170 446116 184226
rect 446184 184170 446240 184226
rect 445812 184046 445868 184102
rect 445936 184046 445992 184102
rect 446060 184046 446116 184102
rect 446184 184046 446240 184102
rect 445812 183922 445868 183978
rect 445936 183922 445992 183978
rect 446060 183922 446116 183978
rect 446184 183922 446240 183978
rect 446612 172294 446668 172350
rect 446736 172294 446792 172350
rect 446860 172294 446916 172350
rect 446984 172294 447040 172350
rect 446612 172170 446668 172226
rect 446736 172170 446792 172226
rect 446860 172170 446916 172226
rect 446984 172170 447040 172226
rect 446612 172046 446668 172102
rect 446736 172046 446792 172102
rect 446860 172046 446916 172102
rect 446984 172046 447040 172102
rect 446612 171922 446668 171978
rect 446736 171922 446792 171978
rect 446860 171922 446916 171978
rect 446984 171922 447040 171978
rect 445812 166294 445868 166350
rect 445936 166294 445992 166350
rect 446060 166294 446116 166350
rect 446184 166294 446240 166350
rect 445812 166170 445868 166226
rect 445936 166170 445992 166226
rect 446060 166170 446116 166226
rect 446184 166170 446240 166226
rect 445812 166046 445868 166102
rect 445936 166046 445992 166102
rect 446060 166046 446116 166102
rect 446184 166046 446240 166102
rect 445812 165922 445868 165978
rect 445936 165922 445992 165978
rect 446060 165922 446116 165978
rect 446184 165922 446240 165978
rect 445564 142262 445620 142318
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 445812 130294 445868 130350
rect 445936 130294 445992 130350
rect 446060 130294 446116 130350
rect 446184 130294 446240 130350
rect 445812 130170 445868 130226
rect 445936 130170 445992 130226
rect 446060 130170 446116 130226
rect 446184 130170 446240 130226
rect 445812 130046 445868 130102
rect 445936 130046 445992 130102
rect 446060 130046 446116 130102
rect 446184 130046 446240 130102
rect 445812 129922 445868 129978
rect 445936 129922 445992 129978
rect 446060 129922 446116 129978
rect 446184 129922 446240 129978
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 446612 118294 446668 118350
rect 446736 118294 446792 118350
rect 446860 118294 446916 118350
rect 446984 118294 447040 118350
rect 446612 118170 446668 118226
rect 446736 118170 446792 118226
rect 446860 118170 446916 118226
rect 446984 118170 447040 118226
rect 446612 118046 446668 118102
rect 446736 118046 446792 118102
rect 446860 118046 446916 118102
rect 446984 118046 447040 118102
rect 446612 117922 446668 117978
rect 446736 117922 446792 117978
rect 446860 117922 446916 117978
rect 446984 117922 447040 117978
rect 445812 112294 445868 112350
rect 445936 112294 445992 112350
rect 446060 112294 446116 112350
rect 446184 112294 446240 112350
rect 445812 112170 445868 112226
rect 445936 112170 445992 112226
rect 446060 112170 446116 112226
rect 446184 112170 446240 112226
rect 445812 112046 445868 112102
rect 445936 112046 445992 112102
rect 446060 112046 446116 112102
rect 446184 112046 446240 112102
rect 445812 111922 445868 111978
rect 445936 111922 445992 111978
rect 446060 111922 446116 111978
rect 446184 111922 446240 111978
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 446612 100294 446668 100350
rect 446736 100294 446792 100350
rect 446860 100294 446916 100350
rect 446984 100294 447040 100350
rect 446612 100170 446668 100226
rect 446736 100170 446792 100226
rect 446860 100170 446916 100226
rect 446984 100170 447040 100226
rect 446612 100046 446668 100102
rect 446736 100046 446792 100102
rect 446860 100046 446916 100102
rect 446984 100046 447040 100102
rect 446612 99922 446668 99978
rect 446736 99922 446792 99978
rect 446860 99922 446916 99978
rect 446984 99922 447040 99978
rect 445812 94294 445868 94350
rect 445936 94294 445992 94350
rect 446060 94294 446116 94350
rect 446184 94294 446240 94350
rect 445812 94170 445868 94226
rect 445936 94170 445992 94226
rect 446060 94170 446116 94226
rect 446184 94170 446240 94226
rect 445812 94046 445868 94102
rect 445936 94046 445992 94102
rect 446060 94046 446116 94102
rect 446184 94046 446240 94102
rect 445812 93922 445868 93978
rect 445936 93922 445992 93978
rect 446060 93922 446116 93978
rect 446184 93922 446240 93978
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 446612 82294 446668 82350
rect 446736 82294 446792 82350
rect 446860 82294 446916 82350
rect 446984 82294 447040 82350
rect 446612 82170 446668 82226
rect 446736 82170 446792 82226
rect 446860 82170 446916 82226
rect 446984 82170 447040 82226
rect 446612 82046 446668 82102
rect 446736 82046 446792 82102
rect 446860 82046 446916 82102
rect 446984 82046 447040 82102
rect 446612 81922 446668 81978
rect 446736 81922 446792 81978
rect 446860 81922 446916 81978
rect 446984 81922 447040 81978
rect 445812 76294 445868 76350
rect 445936 76294 445992 76350
rect 446060 76294 446116 76350
rect 446184 76294 446240 76350
rect 445812 76170 445868 76226
rect 445936 76170 445992 76226
rect 446060 76170 446116 76226
rect 446184 76170 446240 76226
rect 445812 76046 445868 76102
rect 445936 76046 445992 76102
rect 446060 76046 446116 76102
rect 446184 76046 446240 76102
rect 445812 75922 445868 75978
rect 445936 75922 445992 75978
rect 446060 75922 446116 75978
rect 446184 75922 446240 75978
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 446612 64294 446668 64350
rect 446736 64294 446792 64350
rect 446860 64294 446916 64350
rect 446984 64294 447040 64350
rect 446612 64170 446668 64226
rect 446736 64170 446792 64226
rect 446860 64170 446916 64226
rect 446984 64170 447040 64226
rect 446612 64046 446668 64102
rect 446736 64046 446792 64102
rect 446860 64046 446916 64102
rect 446984 64046 447040 64102
rect 446612 63922 446668 63978
rect 446736 63922 446792 63978
rect 446860 63922 446916 63978
rect 446984 63922 447040 63978
rect 445812 58294 445868 58350
rect 445936 58294 445992 58350
rect 446060 58294 446116 58350
rect 446184 58294 446240 58350
rect 445812 58170 445868 58226
rect 445936 58170 445992 58226
rect 446060 58170 446116 58226
rect 446184 58170 446240 58226
rect 445812 58046 445868 58102
rect 445936 58046 445992 58102
rect 446060 58046 446116 58102
rect 446184 58046 446240 58102
rect 445812 57922 445868 57978
rect 445936 57922 445992 57978
rect 446060 57922 446116 57978
rect 446184 57922 446240 57978
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 446612 46294 446668 46350
rect 446736 46294 446792 46350
rect 446860 46294 446916 46350
rect 446984 46294 447040 46350
rect 446612 46170 446668 46226
rect 446736 46170 446792 46226
rect 446860 46170 446916 46226
rect 446984 46170 447040 46226
rect 446612 46046 446668 46102
rect 446736 46046 446792 46102
rect 446860 46046 446916 46102
rect 446984 46046 447040 46102
rect 446612 45922 446668 45978
rect 446736 45922 446792 45978
rect 446860 45922 446916 45978
rect 446984 45922 447040 45978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 457884 367982 457940 368038
rect 454524 366362 454580 366418
rect 454412 364562 454468 364618
rect 452732 358622 452788 358678
rect 452844 356282 452900 356338
rect 456204 361322 456260 361378
rect 456092 353582 456148 353638
rect 457772 350162 457828 350218
rect 461132 248462 461188 248518
rect 464604 235142 464660 235198
rect 466314 418294 466370 418350
rect 466438 418294 466494 418350
rect 466562 418294 466618 418350
rect 466686 418294 466742 418350
rect 466314 418170 466370 418226
rect 466438 418170 466494 418226
rect 466562 418170 466618 418226
rect 466686 418170 466742 418226
rect 466314 418046 466370 418102
rect 466438 418046 466494 418102
rect 466562 418046 466618 418102
rect 466686 418046 466742 418102
rect 466314 417922 466370 417978
rect 466438 417922 466494 417978
rect 466562 417922 466618 417978
rect 466686 417922 466742 417978
rect 470034 514046 470090 514102
rect 470158 514046 470214 514102
rect 470282 514046 470338 514102
rect 470406 514046 470462 514102
rect 470034 513922 470090 513978
rect 470158 513922 470214 513978
rect 470282 513922 470338 513978
rect 470406 513922 470462 513978
rect 489878 514294 489934 514350
rect 490002 514294 490058 514350
rect 489878 514170 489934 514226
rect 490002 514170 490058 514226
rect 489878 514046 489934 514102
rect 490002 514046 490058 514102
rect 489878 513922 489934 513978
rect 490002 513922 490058 513978
rect 520598 514294 520654 514350
rect 520722 514294 520778 514350
rect 520598 514170 520654 514226
rect 520722 514170 520778 514226
rect 520598 514046 520654 514102
rect 520722 514046 520778 514102
rect 520598 513922 520654 513978
rect 520722 513922 520778 513978
rect 474518 508294 474574 508350
rect 474642 508294 474698 508350
rect 474518 508170 474574 508226
rect 474642 508170 474698 508226
rect 474518 508046 474574 508102
rect 474642 508046 474698 508102
rect 474518 507922 474574 507978
rect 474642 507922 474698 507978
rect 505238 508294 505294 508350
rect 505362 508294 505418 508350
rect 505238 508170 505294 508226
rect 505362 508170 505418 508226
rect 505238 508046 505294 508102
rect 505362 508046 505418 508102
rect 505238 507922 505294 507978
rect 505362 507922 505418 507978
rect 535958 508294 536014 508350
rect 536082 508294 536138 508350
rect 535958 508170 536014 508226
rect 536082 508170 536138 508226
rect 535958 508046 536014 508102
rect 536082 508046 536138 508102
rect 535958 507922 536014 507978
rect 536082 507922 536138 507978
rect 470034 496294 470090 496350
rect 470158 496294 470214 496350
rect 470282 496294 470338 496350
rect 470406 496294 470462 496350
rect 470034 496170 470090 496226
rect 470158 496170 470214 496226
rect 470282 496170 470338 496226
rect 470406 496170 470462 496226
rect 470034 496046 470090 496102
rect 470158 496046 470214 496102
rect 470282 496046 470338 496102
rect 470406 496046 470462 496102
rect 470034 495922 470090 495978
rect 470158 495922 470214 495978
rect 470282 495922 470338 495978
rect 470406 495922 470462 495978
rect 474908 499742 474964 499798
rect 474518 490294 474574 490350
rect 474642 490294 474698 490350
rect 474518 490170 474574 490226
rect 474642 490170 474698 490226
rect 474518 490046 474574 490102
rect 474642 490046 474698 490102
rect 474518 489922 474574 489978
rect 474642 489922 474698 489978
rect 470034 478294 470090 478350
rect 470158 478294 470214 478350
rect 470282 478294 470338 478350
rect 470406 478294 470462 478350
rect 470034 478170 470090 478226
rect 470158 478170 470214 478226
rect 470282 478170 470338 478226
rect 470406 478170 470462 478226
rect 470034 478046 470090 478102
rect 470158 478046 470214 478102
rect 470282 478046 470338 478102
rect 470406 478046 470462 478102
rect 470034 477922 470090 477978
rect 470158 477922 470214 477978
rect 470282 477922 470338 477978
rect 470406 477922 470462 477978
rect 474518 472294 474574 472350
rect 474642 472294 474698 472350
rect 474518 472170 474574 472226
rect 474642 472170 474698 472226
rect 474518 472046 474574 472102
rect 474642 472046 474698 472102
rect 474518 471922 474574 471978
rect 474642 471922 474698 471978
rect 470034 460294 470090 460350
rect 470158 460294 470214 460350
rect 470282 460294 470338 460350
rect 470406 460294 470462 460350
rect 470034 460170 470090 460226
rect 470158 460170 470214 460226
rect 470282 460170 470338 460226
rect 470406 460170 470462 460226
rect 470034 460046 470090 460102
rect 470158 460046 470214 460102
rect 470282 460046 470338 460102
rect 470406 460046 470462 460102
rect 470034 459922 470090 459978
rect 470158 459922 470214 459978
rect 470282 459922 470338 459978
rect 470406 459922 470462 459978
rect 474518 454294 474574 454350
rect 474642 454294 474698 454350
rect 474518 454170 474574 454226
rect 474642 454170 474698 454226
rect 474518 454046 474574 454102
rect 474642 454046 474698 454102
rect 474518 453922 474574 453978
rect 474642 453922 474698 453978
rect 489878 496294 489934 496350
rect 490002 496294 490058 496350
rect 489878 496170 489934 496226
rect 490002 496170 490058 496226
rect 489878 496046 489934 496102
rect 490002 496046 490058 496102
rect 489878 495922 489934 495978
rect 490002 495922 490058 495978
rect 520598 496294 520654 496350
rect 520722 496294 520778 496350
rect 520598 496170 520654 496226
rect 520722 496170 520778 496226
rect 520598 496046 520654 496102
rect 520722 496046 520778 496102
rect 520598 495922 520654 495978
rect 520722 495922 520778 495978
rect 505238 490294 505294 490350
rect 505362 490294 505418 490350
rect 505238 490170 505294 490226
rect 505362 490170 505418 490226
rect 505238 490046 505294 490102
rect 505362 490046 505418 490102
rect 505238 489922 505294 489978
rect 505362 489922 505418 489978
rect 535958 490294 536014 490350
rect 536082 490294 536138 490350
rect 535958 490170 536014 490226
rect 536082 490170 536138 490226
rect 535958 490046 536014 490102
rect 536082 490046 536138 490102
rect 535958 489922 536014 489978
rect 536082 489922 536138 489978
rect 489878 478294 489934 478350
rect 490002 478294 490058 478350
rect 489878 478170 489934 478226
rect 490002 478170 490058 478226
rect 489878 478046 489934 478102
rect 490002 478046 490058 478102
rect 489878 477922 489934 477978
rect 490002 477922 490058 477978
rect 520598 478294 520654 478350
rect 520722 478294 520778 478350
rect 520598 478170 520654 478226
rect 520722 478170 520778 478226
rect 520598 478046 520654 478102
rect 520722 478046 520778 478102
rect 520598 477922 520654 477978
rect 520722 477922 520778 477978
rect 505238 472294 505294 472350
rect 505362 472294 505418 472350
rect 505238 472170 505294 472226
rect 505362 472170 505418 472226
rect 505238 472046 505294 472102
rect 505362 472046 505418 472102
rect 505238 471922 505294 471978
rect 505362 471922 505418 471978
rect 535958 472294 536014 472350
rect 536082 472294 536138 472350
rect 535958 472170 536014 472226
rect 536082 472170 536138 472226
rect 535958 472046 536014 472102
rect 536082 472046 536138 472102
rect 535958 471922 536014 471978
rect 536082 471922 536138 471978
rect 489878 460294 489934 460350
rect 490002 460294 490058 460350
rect 489878 460170 489934 460226
rect 490002 460170 490058 460226
rect 489878 460046 489934 460102
rect 490002 460046 490058 460102
rect 489878 459922 489934 459978
rect 490002 459922 490058 459978
rect 520598 460294 520654 460350
rect 520722 460294 520778 460350
rect 520598 460170 520654 460226
rect 520722 460170 520778 460226
rect 520598 460046 520654 460102
rect 520722 460046 520778 460102
rect 520598 459922 520654 459978
rect 520722 459922 520778 459978
rect 505238 454294 505294 454350
rect 505362 454294 505418 454350
rect 505238 454170 505294 454226
rect 505362 454170 505418 454226
rect 505238 454046 505294 454102
rect 505362 454046 505418 454102
rect 505238 453922 505294 453978
rect 505362 453922 505418 453978
rect 535958 454294 536014 454350
rect 536082 454294 536138 454350
rect 535958 454170 536014 454226
rect 536082 454170 536138 454226
rect 535958 454046 536014 454102
rect 536082 454046 536138 454102
rect 535958 453922 536014 453978
rect 536082 453922 536138 453978
rect 478044 450962 478100 451018
rect 470034 442294 470090 442350
rect 470158 442294 470214 442350
rect 470282 442294 470338 442350
rect 470406 442294 470462 442350
rect 470034 442170 470090 442226
rect 470158 442170 470214 442226
rect 470282 442170 470338 442226
rect 470406 442170 470462 442226
rect 470034 442046 470090 442102
rect 470158 442046 470214 442102
rect 470282 442046 470338 442102
rect 470406 442046 470462 442102
rect 470034 441922 470090 441978
rect 470158 441922 470214 441978
rect 470282 441922 470338 441978
rect 470406 441922 470462 441978
rect 470034 424294 470090 424350
rect 470158 424294 470214 424350
rect 470282 424294 470338 424350
rect 470406 424294 470462 424350
rect 470034 424170 470090 424226
rect 470158 424170 470214 424226
rect 470282 424170 470338 424226
rect 470406 424170 470462 424226
rect 470034 424046 470090 424102
rect 470158 424046 470214 424102
rect 470282 424046 470338 424102
rect 470406 424046 470462 424102
rect 470034 423922 470090 423978
rect 470158 423922 470214 423978
rect 470282 423922 470338 423978
rect 470406 423922 470462 423978
rect 470034 406294 470090 406350
rect 470158 406294 470214 406350
rect 470282 406294 470338 406350
rect 470406 406294 470462 406350
rect 470034 406170 470090 406226
rect 470158 406170 470214 406226
rect 470282 406170 470338 406226
rect 470406 406170 470462 406226
rect 470034 406046 470090 406102
rect 470158 406046 470214 406102
rect 470282 406046 470338 406102
rect 470406 406046 470462 406102
rect 470034 405922 470090 405978
rect 470158 405922 470214 405978
rect 470282 405922 470338 405978
rect 470406 405922 470462 405978
rect 467852 404342 467908 404398
rect 468636 404342 468692 404398
rect 466314 400294 466370 400350
rect 466438 400294 466494 400350
rect 466562 400294 466618 400350
rect 466686 400294 466742 400350
rect 466314 400170 466370 400226
rect 466438 400170 466494 400226
rect 466562 400170 466618 400226
rect 466686 400170 466742 400226
rect 466314 400046 466370 400102
rect 466438 400046 466494 400102
rect 466562 400046 466618 400102
rect 466686 400046 466742 400102
rect 466314 399922 466370 399978
rect 466438 399922 466494 399978
rect 466562 399922 466618 399978
rect 466686 399922 466742 399978
rect 466314 382294 466370 382350
rect 466438 382294 466494 382350
rect 466562 382294 466618 382350
rect 466686 382294 466742 382350
rect 466314 382170 466370 382226
rect 466438 382170 466494 382226
rect 466562 382170 466618 382226
rect 466686 382170 466742 382226
rect 466314 382046 466370 382102
rect 466438 382046 466494 382102
rect 466562 382046 466618 382102
rect 466686 382046 466742 382102
rect 466314 381922 466370 381978
rect 466438 381922 466494 381978
rect 466562 381922 466618 381978
rect 466686 381922 466742 381978
rect 466314 364294 466370 364350
rect 466438 364294 466494 364350
rect 466562 364294 466618 364350
rect 466686 364294 466742 364350
rect 466314 364170 466370 364226
rect 466438 364170 466494 364226
rect 466562 364170 466618 364226
rect 466686 364170 466742 364226
rect 466314 364046 466370 364102
rect 466438 364046 466494 364102
rect 466562 364046 466618 364102
rect 466686 364046 466742 364102
rect 466314 363922 466370 363978
rect 466438 363922 466494 363978
rect 466562 363922 466618 363978
rect 466686 363922 466742 363978
rect 466314 346294 466370 346350
rect 466438 346294 466494 346350
rect 466562 346294 466618 346350
rect 466686 346294 466742 346350
rect 466314 346170 466370 346226
rect 466438 346170 466494 346226
rect 466562 346170 466618 346226
rect 466686 346170 466742 346226
rect 466314 346046 466370 346102
rect 466438 346046 466494 346102
rect 466562 346046 466618 346102
rect 466686 346046 466742 346102
rect 466314 345922 466370 345978
rect 466438 345922 466494 345978
rect 466562 345922 466618 345978
rect 466686 345922 466742 345978
rect 466314 328294 466370 328350
rect 466438 328294 466494 328350
rect 466562 328294 466618 328350
rect 466686 328294 466742 328350
rect 466314 328170 466370 328226
rect 466438 328170 466494 328226
rect 466562 328170 466618 328226
rect 466686 328170 466742 328226
rect 466314 328046 466370 328102
rect 466438 328046 466494 328102
rect 466562 328046 466618 328102
rect 466686 328046 466742 328102
rect 466314 327922 466370 327978
rect 466438 327922 466494 327978
rect 466562 327922 466618 327978
rect 466686 327922 466742 327978
rect 466314 310294 466370 310350
rect 466438 310294 466494 310350
rect 466562 310294 466618 310350
rect 466686 310294 466742 310350
rect 466314 310170 466370 310226
rect 466438 310170 466494 310226
rect 466562 310170 466618 310226
rect 466686 310170 466742 310226
rect 466314 310046 466370 310102
rect 466438 310046 466494 310102
rect 466562 310046 466618 310102
rect 466686 310046 466742 310102
rect 466314 309922 466370 309978
rect 466438 309922 466494 309978
rect 466562 309922 466618 309978
rect 466686 309922 466742 309978
rect 466314 292294 466370 292350
rect 466438 292294 466494 292350
rect 466562 292294 466618 292350
rect 466686 292294 466742 292350
rect 466314 292170 466370 292226
rect 466438 292170 466494 292226
rect 466562 292170 466618 292226
rect 466686 292170 466742 292226
rect 466314 292046 466370 292102
rect 466438 292046 466494 292102
rect 466562 292046 466618 292102
rect 466686 292046 466742 292102
rect 466314 291922 466370 291978
rect 466438 291922 466494 291978
rect 466562 291922 466618 291978
rect 466686 291922 466742 291978
rect 466314 274294 466370 274350
rect 466438 274294 466494 274350
rect 466562 274294 466618 274350
rect 466686 274294 466742 274350
rect 466314 274170 466370 274226
rect 466438 274170 466494 274226
rect 466562 274170 466618 274226
rect 466686 274170 466742 274226
rect 466314 274046 466370 274102
rect 466438 274046 466494 274102
rect 466562 274046 466618 274102
rect 466686 274046 466742 274102
rect 466314 273922 466370 273978
rect 466438 273922 466494 273978
rect 466562 273922 466618 273978
rect 466686 273922 466742 273978
rect 466314 256294 466370 256350
rect 466438 256294 466494 256350
rect 466562 256294 466618 256350
rect 466686 256294 466742 256350
rect 466314 256170 466370 256226
rect 466438 256170 466494 256226
rect 466562 256170 466618 256226
rect 466686 256170 466742 256226
rect 466314 256046 466370 256102
rect 466438 256046 466494 256102
rect 466562 256046 466618 256102
rect 466686 256046 466742 256102
rect 466314 255922 466370 255978
rect 466438 255922 466494 255978
rect 466562 255922 466618 255978
rect 466686 255922 466742 255978
rect 466314 238294 466370 238350
rect 466438 238294 466494 238350
rect 466562 238294 466618 238350
rect 466686 238294 466742 238350
rect 466314 238170 466370 238226
rect 466438 238170 466494 238226
rect 466562 238170 466618 238226
rect 466686 238170 466742 238226
rect 466314 238046 466370 238102
rect 466438 238046 466494 238102
rect 466562 238046 466618 238102
rect 466686 238046 466742 238102
rect 466314 237922 466370 237978
rect 466438 237922 466494 237978
rect 466562 237922 466618 237978
rect 466686 237922 466742 237978
rect 464492 206522 464548 206578
rect 466314 220294 466370 220350
rect 466438 220294 466494 220350
rect 466562 220294 466618 220350
rect 466686 220294 466742 220350
rect 466314 220170 466370 220226
rect 466438 220170 466494 220226
rect 466562 220170 466618 220226
rect 466686 220170 466742 220226
rect 466314 220046 466370 220102
rect 466438 220046 466494 220102
rect 466562 220046 466618 220102
rect 466686 220046 466742 220102
rect 466314 219922 466370 219978
rect 466438 219922 466494 219978
rect 466562 219922 466618 219978
rect 466686 219922 466742 219978
rect 466314 202294 466370 202350
rect 466438 202294 466494 202350
rect 466562 202294 466618 202350
rect 466686 202294 466742 202350
rect 466314 202170 466370 202226
rect 466438 202170 466494 202226
rect 466562 202170 466618 202226
rect 466686 202170 466742 202226
rect 466314 202046 466370 202102
rect 466438 202046 466494 202102
rect 466562 202046 466618 202102
rect 466686 202046 466742 202102
rect 466314 201922 466370 201978
rect 466438 201922 466494 201978
rect 466562 201922 466618 201978
rect 466686 201922 466742 201978
rect 466314 184294 466370 184350
rect 466438 184294 466494 184350
rect 466562 184294 466618 184350
rect 466686 184294 466742 184350
rect 466314 184170 466370 184226
rect 466438 184170 466494 184226
rect 466562 184170 466618 184226
rect 466686 184170 466742 184226
rect 466314 184046 466370 184102
rect 466438 184046 466494 184102
rect 466562 184046 466618 184102
rect 466686 184046 466742 184102
rect 466314 183922 466370 183978
rect 466438 183922 466494 183978
rect 466562 183922 466618 183978
rect 466686 183922 466742 183978
rect 466314 166294 466370 166350
rect 466438 166294 466494 166350
rect 466562 166294 466618 166350
rect 466686 166294 466742 166350
rect 466314 166170 466370 166226
rect 466438 166170 466494 166226
rect 466562 166170 466618 166226
rect 466686 166170 466742 166226
rect 466314 166046 466370 166102
rect 466438 166046 466494 166102
rect 466562 166046 466618 166102
rect 466686 166046 466742 166102
rect 466314 165922 466370 165978
rect 466438 165922 466494 165978
rect 466562 165922 466618 165978
rect 466686 165922 466742 165978
rect 466314 148294 466370 148350
rect 466438 148294 466494 148350
rect 466562 148294 466618 148350
rect 466686 148294 466742 148350
rect 466314 148170 466370 148226
rect 466438 148170 466494 148226
rect 466562 148170 466618 148226
rect 466686 148170 466742 148226
rect 466314 148046 466370 148102
rect 466438 148046 466494 148102
rect 466562 148046 466618 148102
rect 466686 148046 466742 148102
rect 466314 147922 466370 147978
rect 466438 147922 466494 147978
rect 466562 147922 466618 147978
rect 466686 147922 466742 147978
rect 461130 130294 461186 130350
rect 461254 130294 461310 130350
rect 461378 130294 461434 130350
rect 461502 130294 461558 130350
rect 461130 130170 461186 130226
rect 461254 130170 461310 130226
rect 461378 130170 461434 130226
rect 461502 130170 461558 130226
rect 461130 130046 461186 130102
rect 461254 130046 461310 130102
rect 461378 130046 461434 130102
rect 461502 130046 461558 130102
rect 461130 129922 461186 129978
rect 461254 129922 461310 129978
rect 461378 129922 461434 129978
rect 461502 129922 461558 129978
rect 466314 130294 466370 130350
rect 466438 130294 466494 130350
rect 466562 130294 466618 130350
rect 466686 130294 466742 130350
rect 466314 130170 466370 130226
rect 466438 130170 466494 130226
rect 466562 130170 466618 130226
rect 466686 130170 466742 130226
rect 466314 130046 466370 130102
rect 466438 130046 466494 130102
rect 466562 130046 466618 130102
rect 466686 130046 466742 130102
rect 466314 129922 466370 129978
rect 466438 129922 466494 129978
rect 466562 129922 466618 129978
rect 466686 129922 466742 129978
rect 461930 118294 461986 118350
rect 462054 118294 462110 118350
rect 462178 118294 462234 118350
rect 462302 118294 462358 118350
rect 461930 118170 461986 118226
rect 462054 118170 462110 118226
rect 462178 118170 462234 118226
rect 462302 118170 462358 118226
rect 461930 118046 461986 118102
rect 462054 118046 462110 118102
rect 462178 118046 462234 118102
rect 462302 118046 462358 118102
rect 461930 117922 461986 117978
rect 462054 117922 462110 117978
rect 462178 117922 462234 117978
rect 462302 117922 462358 117978
rect 461130 112294 461186 112350
rect 461254 112294 461310 112350
rect 461378 112294 461434 112350
rect 461502 112294 461558 112350
rect 461130 112170 461186 112226
rect 461254 112170 461310 112226
rect 461378 112170 461434 112226
rect 461502 112170 461558 112226
rect 461130 112046 461186 112102
rect 461254 112046 461310 112102
rect 461378 112046 461434 112102
rect 461502 112046 461558 112102
rect 461130 111922 461186 111978
rect 461254 111922 461310 111978
rect 461378 111922 461434 111978
rect 461502 111922 461558 111978
rect 466314 112294 466370 112350
rect 466438 112294 466494 112350
rect 466562 112294 466618 112350
rect 466686 112294 466742 112350
rect 466314 112170 466370 112226
rect 466438 112170 466494 112226
rect 466562 112170 466618 112226
rect 466686 112170 466742 112226
rect 466314 112046 466370 112102
rect 466438 112046 466494 112102
rect 466562 112046 466618 112102
rect 466686 112046 466742 112102
rect 466314 111922 466370 111978
rect 466438 111922 466494 111978
rect 466562 111922 466618 111978
rect 466686 111922 466742 111978
rect 461930 100294 461986 100350
rect 462054 100294 462110 100350
rect 462178 100294 462234 100350
rect 462302 100294 462358 100350
rect 461930 100170 461986 100226
rect 462054 100170 462110 100226
rect 462178 100170 462234 100226
rect 462302 100170 462358 100226
rect 461930 100046 461986 100102
rect 462054 100046 462110 100102
rect 462178 100046 462234 100102
rect 462302 100046 462358 100102
rect 461930 99922 461986 99978
rect 462054 99922 462110 99978
rect 462178 99922 462234 99978
rect 462302 99922 462358 99978
rect 461130 94294 461186 94350
rect 461254 94294 461310 94350
rect 461378 94294 461434 94350
rect 461502 94294 461558 94350
rect 461130 94170 461186 94226
rect 461254 94170 461310 94226
rect 461378 94170 461434 94226
rect 461502 94170 461558 94226
rect 461130 94046 461186 94102
rect 461254 94046 461310 94102
rect 461378 94046 461434 94102
rect 461502 94046 461558 94102
rect 461130 93922 461186 93978
rect 461254 93922 461310 93978
rect 461378 93922 461434 93978
rect 461502 93922 461558 93978
rect 466314 94294 466370 94350
rect 466438 94294 466494 94350
rect 466562 94294 466618 94350
rect 466686 94294 466742 94350
rect 466314 94170 466370 94226
rect 466438 94170 466494 94226
rect 466562 94170 466618 94226
rect 466686 94170 466742 94226
rect 466314 94046 466370 94102
rect 466438 94046 466494 94102
rect 466562 94046 466618 94102
rect 466686 94046 466742 94102
rect 466314 93922 466370 93978
rect 466438 93922 466494 93978
rect 466562 93922 466618 93978
rect 466686 93922 466742 93978
rect 461930 82294 461986 82350
rect 462054 82294 462110 82350
rect 462178 82294 462234 82350
rect 462302 82294 462358 82350
rect 461930 82170 461986 82226
rect 462054 82170 462110 82226
rect 462178 82170 462234 82226
rect 462302 82170 462358 82226
rect 461930 82046 461986 82102
rect 462054 82046 462110 82102
rect 462178 82046 462234 82102
rect 462302 82046 462358 82102
rect 461930 81922 461986 81978
rect 462054 81922 462110 81978
rect 462178 81922 462234 81978
rect 462302 81922 462358 81978
rect 461130 76294 461186 76350
rect 461254 76294 461310 76350
rect 461378 76294 461434 76350
rect 461502 76294 461558 76350
rect 461130 76170 461186 76226
rect 461254 76170 461310 76226
rect 461378 76170 461434 76226
rect 461502 76170 461558 76226
rect 461130 76046 461186 76102
rect 461254 76046 461310 76102
rect 461378 76046 461434 76102
rect 461502 76046 461558 76102
rect 461130 75922 461186 75978
rect 461254 75922 461310 75978
rect 461378 75922 461434 75978
rect 461502 75922 461558 75978
rect 466314 76294 466370 76350
rect 466438 76294 466494 76350
rect 466562 76294 466618 76350
rect 466686 76294 466742 76350
rect 466314 76170 466370 76226
rect 466438 76170 466494 76226
rect 466562 76170 466618 76226
rect 466686 76170 466742 76226
rect 466314 76046 466370 76102
rect 466438 76046 466494 76102
rect 466562 76046 466618 76102
rect 466686 76046 466742 76102
rect 466314 75922 466370 75978
rect 466438 75922 466494 75978
rect 466562 75922 466618 75978
rect 466686 75922 466742 75978
rect 461930 64294 461986 64350
rect 462054 64294 462110 64350
rect 462178 64294 462234 64350
rect 462302 64294 462358 64350
rect 461930 64170 461986 64226
rect 462054 64170 462110 64226
rect 462178 64170 462234 64226
rect 462302 64170 462358 64226
rect 461930 64046 461986 64102
rect 462054 64046 462110 64102
rect 462178 64046 462234 64102
rect 462302 64046 462358 64102
rect 461930 63922 461986 63978
rect 462054 63922 462110 63978
rect 462178 63922 462234 63978
rect 462302 63922 462358 63978
rect 461130 58294 461186 58350
rect 461254 58294 461310 58350
rect 461378 58294 461434 58350
rect 461502 58294 461558 58350
rect 461130 58170 461186 58226
rect 461254 58170 461310 58226
rect 461378 58170 461434 58226
rect 461502 58170 461558 58226
rect 461130 58046 461186 58102
rect 461254 58046 461310 58102
rect 461378 58046 461434 58102
rect 461502 58046 461558 58102
rect 461130 57922 461186 57978
rect 461254 57922 461310 57978
rect 461378 57922 461434 57978
rect 461502 57922 461558 57978
rect 466314 58294 466370 58350
rect 466438 58294 466494 58350
rect 466562 58294 466618 58350
rect 466686 58294 466742 58350
rect 466314 58170 466370 58226
rect 466438 58170 466494 58226
rect 466562 58170 466618 58226
rect 466686 58170 466742 58226
rect 466314 58046 466370 58102
rect 466438 58046 466494 58102
rect 466562 58046 466618 58102
rect 466686 58046 466742 58102
rect 466314 57922 466370 57978
rect 466438 57922 466494 57978
rect 466562 57922 466618 57978
rect 466686 57922 466742 57978
rect 461930 46294 461986 46350
rect 462054 46294 462110 46350
rect 462178 46294 462234 46350
rect 462302 46294 462358 46350
rect 461930 46170 461986 46226
rect 462054 46170 462110 46226
rect 462178 46170 462234 46226
rect 462302 46170 462358 46226
rect 461930 46046 461986 46102
rect 462054 46046 462110 46102
rect 462178 46046 462234 46102
rect 462302 46046 462358 46102
rect 461930 45922 461986 45978
rect 462054 45922 462110 45978
rect 462178 45922 462234 45978
rect 462302 45922 462358 45978
rect 466314 40294 466370 40350
rect 466438 40294 466494 40350
rect 466562 40294 466618 40350
rect 466686 40294 466742 40350
rect 466314 40170 466370 40226
rect 466438 40170 466494 40226
rect 466562 40170 466618 40226
rect 466686 40170 466742 40226
rect 466314 40046 466370 40102
rect 466438 40046 466494 40102
rect 466562 40046 466618 40102
rect 466686 40046 466742 40102
rect 466314 39922 466370 39978
rect 466438 39922 466494 39978
rect 466562 39922 466618 39978
rect 466686 39922 466742 39978
rect 466314 22294 466370 22350
rect 466438 22294 466494 22350
rect 466562 22294 466618 22350
rect 466686 22294 466742 22350
rect 466314 22170 466370 22226
rect 466438 22170 466494 22226
rect 466562 22170 466618 22226
rect 466686 22170 466742 22226
rect 466314 22046 466370 22102
rect 466438 22046 466494 22102
rect 466562 22046 466618 22102
rect 466686 22046 466742 22102
rect 466314 21922 466370 21978
rect 466438 21922 466494 21978
rect 466562 21922 466618 21978
rect 466686 21922 466742 21978
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 470034 388294 470090 388350
rect 470158 388294 470214 388350
rect 470282 388294 470338 388350
rect 470406 388294 470462 388350
rect 470034 388170 470090 388226
rect 470158 388170 470214 388226
rect 470282 388170 470338 388226
rect 470406 388170 470462 388226
rect 470034 388046 470090 388102
rect 470158 388046 470214 388102
rect 470282 388046 470338 388102
rect 470406 388046 470462 388102
rect 470034 387922 470090 387978
rect 470158 387922 470214 387978
rect 470282 387922 470338 387978
rect 470406 387922 470462 387978
rect 470034 370294 470090 370350
rect 470158 370294 470214 370350
rect 470282 370294 470338 370350
rect 470406 370294 470462 370350
rect 470034 370170 470090 370226
rect 470158 370170 470214 370226
rect 470282 370170 470338 370226
rect 470406 370170 470462 370226
rect 470034 370046 470090 370102
rect 470158 370046 470214 370102
rect 470282 370046 470338 370102
rect 470406 370046 470462 370102
rect 470034 369922 470090 369978
rect 470158 369922 470214 369978
rect 470282 369922 470338 369978
rect 470406 369922 470462 369978
rect 470034 352294 470090 352350
rect 470158 352294 470214 352350
rect 470282 352294 470338 352350
rect 470406 352294 470462 352350
rect 470034 352170 470090 352226
rect 470158 352170 470214 352226
rect 470282 352170 470338 352226
rect 470406 352170 470462 352226
rect 470034 352046 470090 352102
rect 470158 352046 470214 352102
rect 470282 352046 470338 352102
rect 470406 352046 470462 352102
rect 470034 351922 470090 351978
rect 470158 351922 470214 351978
rect 470282 351922 470338 351978
rect 470406 351922 470462 351978
rect 470034 334294 470090 334350
rect 470158 334294 470214 334350
rect 470282 334294 470338 334350
rect 470406 334294 470462 334350
rect 470034 334170 470090 334226
rect 470158 334170 470214 334226
rect 470282 334170 470338 334226
rect 470406 334170 470462 334226
rect 470034 334046 470090 334102
rect 470158 334046 470214 334102
rect 470282 334046 470338 334102
rect 470406 334046 470462 334102
rect 470034 333922 470090 333978
rect 470158 333922 470214 333978
rect 470282 333922 470338 333978
rect 470406 333922 470462 333978
rect 470034 316294 470090 316350
rect 470158 316294 470214 316350
rect 470282 316294 470338 316350
rect 470406 316294 470462 316350
rect 470034 316170 470090 316226
rect 470158 316170 470214 316226
rect 470282 316170 470338 316226
rect 470406 316170 470462 316226
rect 470034 316046 470090 316102
rect 470158 316046 470214 316102
rect 470282 316046 470338 316102
rect 470406 316046 470462 316102
rect 470034 315922 470090 315978
rect 470158 315922 470214 315978
rect 470282 315922 470338 315978
rect 470406 315922 470462 315978
rect 470034 298294 470090 298350
rect 470158 298294 470214 298350
rect 470282 298294 470338 298350
rect 470406 298294 470462 298350
rect 470034 298170 470090 298226
rect 470158 298170 470214 298226
rect 470282 298170 470338 298226
rect 470406 298170 470462 298226
rect 470034 298046 470090 298102
rect 470158 298046 470214 298102
rect 470282 298046 470338 298102
rect 470406 298046 470462 298102
rect 470034 297922 470090 297978
rect 470158 297922 470214 297978
rect 470282 297922 470338 297978
rect 470406 297922 470462 297978
rect 477932 431882 477988 431938
rect 475692 340262 475748 340318
rect 475468 339182 475524 339238
rect 475468 337562 475524 337618
rect 475580 337382 475636 337438
rect 475468 335942 475524 335998
rect 475468 333602 475524 333658
rect 475468 332522 475524 332578
rect 475580 332342 475636 332398
rect 475468 330902 475524 330958
rect 476252 340082 476308 340138
rect 475468 326042 475524 326098
rect 475468 321002 475524 321058
rect 475468 317772 475524 317818
rect 475468 317762 475524 317772
rect 475580 317582 475636 317638
rect 475468 314162 475524 314218
rect 475468 312542 475524 312598
rect 475468 307502 475524 307558
rect 474572 300482 474628 300538
rect 476140 290582 476196 290638
rect 476028 288422 476084 288478
rect 475468 283562 475524 283618
rect 476364 285362 476420 285418
rect 476700 290402 476756 290458
rect 476588 287162 476644 287218
rect 476924 293642 476980 293698
rect 476812 286982 476868 287038
rect 477036 286802 477092 286858
rect 470034 280294 470090 280350
rect 470158 280294 470214 280350
rect 470282 280294 470338 280350
rect 470406 280294 470462 280350
rect 470034 280170 470090 280226
rect 470158 280170 470214 280226
rect 470282 280170 470338 280226
rect 470406 280170 470462 280226
rect 470034 280046 470090 280102
rect 470158 280046 470214 280102
rect 470282 280046 470338 280102
rect 470406 280046 470462 280102
rect 470034 279922 470090 279978
rect 470158 279922 470214 279978
rect 470282 279922 470338 279978
rect 470406 279922 470462 279978
rect 479836 432422 479892 432478
rect 478492 404522 478548 404578
rect 479612 432242 479668 432298
rect 478156 288602 478212 288658
rect 479724 295082 479780 295138
rect 480060 432062 480116 432118
rect 479948 295262 480004 295318
rect 480620 405422 480676 405478
rect 512316 433322 512372 433378
rect 498876 432422 498932 432478
rect 481628 405422 481684 405478
rect 481516 403082 481572 403138
rect 481404 402902 481460 402958
rect 502908 432242 502964 432298
rect 519036 432062 519092 432118
rect 499878 424294 499934 424350
rect 500002 424294 500058 424350
rect 499878 424170 499934 424226
rect 500002 424170 500058 424226
rect 499878 424046 499934 424102
rect 500002 424046 500058 424102
rect 499878 423922 499934 423978
rect 500002 423922 500058 423978
rect 484518 418294 484574 418350
rect 484642 418294 484698 418350
rect 484518 418170 484574 418226
rect 484642 418170 484698 418226
rect 484518 418046 484574 418102
rect 484642 418046 484698 418102
rect 484518 417922 484574 417978
rect 484642 417922 484698 417978
rect 515238 418294 515294 418350
rect 515362 418294 515418 418350
rect 515238 418170 515294 418226
rect 515362 418170 515418 418226
rect 515238 418046 515294 418102
rect 515362 418046 515418 418102
rect 515238 417922 515294 417978
rect 515362 417922 515418 417978
rect 499878 406294 499934 406350
rect 500002 406294 500058 406350
rect 499878 406170 499934 406226
rect 500002 406170 500058 406226
rect 499878 406046 499934 406102
rect 500002 406046 500058 406102
rect 499878 405922 499934 405978
rect 500002 405922 500058 405978
rect 483084 402722 483140 402778
rect 484518 400294 484574 400350
rect 484642 400294 484698 400350
rect 484518 400170 484574 400226
rect 484642 400170 484698 400226
rect 484518 400046 484574 400102
rect 484642 400046 484698 400102
rect 484518 399922 484574 399978
rect 484642 399922 484698 399978
rect 515238 400294 515294 400350
rect 515362 400294 515418 400350
rect 515238 400170 515294 400226
rect 515362 400170 515418 400226
rect 515238 400046 515294 400102
rect 515362 400046 515418 400102
rect 515238 399922 515294 399978
rect 515362 399922 515418 399978
rect 482972 398042 483028 398098
rect 499878 388294 499934 388350
rect 500002 388294 500058 388350
rect 499878 388170 499934 388226
rect 500002 388170 500058 388226
rect 499878 388046 499934 388102
rect 500002 388046 500058 388102
rect 499878 387922 499934 387978
rect 500002 387922 500058 387978
rect 497034 382294 497090 382350
rect 497158 382294 497214 382350
rect 497282 382294 497338 382350
rect 497406 382294 497462 382350
rect 497034 382170 497090 382226
rect 497158 382170 497214 382226
rect 497282 382170 497338 382226
rect 497406 382170 497462 382226
rect 497034 382046 497090 382102
rect 497158 382046 497214 382102
rect 497282 382046 497338 382102
rect 497406 382046 497462 382102
rect 497034 381922 497090 381978
rect 497158 381922 497214 381978
rect 497282 381922 497338 381978
rect 497406 381922 497462 381978
rect 494844 377702 494900 377758
rect 498876 377522 498932 377578
rect 497034 364294 497090 364350
rect 497158 364294 497214 364350
rect 497282 364294 497338 364350
rect 497406 364294 497462 364350
rect 497034 364170 497090 364226
rect 497158 364170 497214 364226
rect 497282 364170 497338 364226
rect 497406 364170 497462 364226
rect 497034 364046 497090 364102
rect 497158 364046 497214 364102
rect 497282 364046 497338 364102
rect 497406 364046 497462 364102
rect 497034 363922 497090 363978
rect 497158 363922 497214 363978
rect 497282 363922 497338 363978
rect 497406 363922 497462 363978
rect 495964 348542 496020 348598
rect 521052 377916 521108 377938
rect 521052 377882 521108 377916
rect 523068 431882 523124 431938
rect 525868 388862 525924 388918
rect 526652 388862 526708 388918
rect 527754 436294 527810 436350
rect 527878 436294 527934 436350
rect 528002 436294 528058 436350
rect 528126 436294 528182 436350
rect 527754 436170 527810 436226
rect 527878 436170 527934 436226
rect 528002 436170 528058 436226
rect 528126 436170 528182 436226
rect 527754 436046 527810 436102
rect 527878 436046 527934 436102
rect 528002 436046 528058 436102
rect 528126 436046 528182 436102
rect 527754 435922 527810 435978
rect 527878 435922 527934 435978
rect 528002 435922 528058 435978
rect 528126 435922 528182 435978
rect 527754 418294 527810 418350
rect 527878 418294 527934 418350
rect 528002 418294 528058 418350
rect 528126 418294 528182 418350
rect 527754 418170 527810 418226
rect 527878 418170 527934 418226
rect 528002 418170 528058 418226
rect 528126 418170 528182 418226
rect 527754 418046 527810 418102
rect 527878 418046 527934 418102
rect 528002 418046 528058 418102
rect 528126 418046 528182 418102
rect 527754 417922 527810 417978
rect 527878 417922 527934 417978
rect 528002 417922 528058 417978
rect 528126 417922 528182 417978
rect 527754 400294 527810 400350
rect 527878 400294 527934 400350
rect 528002 400294 528058 400350
rect 528126 400294 528182 400350
rect 527754 400170 527810 400226
rect 527878 400170 527934 400226
rect 528002 400170 528058 400226
rect 528126 400170 528182 400226
rect 527754 400046 527810 400102
rect 527878 400046 527934 400102
rect 528002 400046 528058 400102
rect 528126 400046 528182 400102
rect 527754 399922 527810 399978
rect 527878 399922 527934 399978
rect 528002 399922 528058 399978
rect 528126 399922 528182 399978
rect 527754 382294 527810 382350
rect 527878 382294 527934 382350
rect 528002 382294 528058 382350
rect 528126 382294 528182 382350
rect 527754 382170 527810 382226
rect 527878 382170 527934 382226
rect 528002 382170 528058 382226
rect 528126 382170 528182 382226
rect 527754 382046 527810 382102
rect 527878 382046 527934 382102
rect 528002 382046 528058 382102
rect 528126 382046 528182 382102
rect 527754 381922 527810 381978
rect 527878 381922 527934 381978
rect 528002 381922 528058 381978
rect 528126 381922 528182 381978
rect 500754 370294 500810 370350
rect 500878 370294 500934 370350
rect 501002 370294 501058 370350
rect 501126 370294 501182 370350
rect 500754 370170 500810 370226
rect 500878 370170 500934 370226
rect 501002 370170 501058 370226
rect 501126 370170 501182 370226
rect 500754 370046 500810 370102
rect 500878 370046 500934 370102
rect 501002 370046 501058 370102
rect 501126 370046 501182 370102
rect 500754 369922 500810 369978
rect 500878 369922 500934 369978
rect 501002 369922 501058 369978
rect 501126 369922 501182 369978
rect 497034 346294 497090 346350
rect 497158 346294 497214 346350
rect 497282 346294 497338 346350
rect 497406 346294 497462 346350
rect 497034 346170 497090 346226
rect 497158 346170 497214 346226
rect 497282 346170 497338 346226
rect 497406 346170 497462 346226
rect 497034 346046 497090 346102
rect 497158 346046 497214 346102
rect 497282 346046 497338 346102
rect 497406 346046 497462 346102
rect 497034 345922 497090 345978
rect 497158 345922 497214 345978
rect 497282 345922 497338 345978
rect 497406 345922 497462 345978
rect 498988 360242 499044 360298
rect 505708 373742 505764 373798
rect 500754 352294 500810 352350
rect 500878 352294 500934 352350
rect 501002 352294 501058 352350
rect 501126 352294 501182 352350
rect 500754 352170 500810 352226
rect 500878 352170 500934 352226
rect 501002 352170 501058 352226
rect 501126 352170 501182 352226
rect 500754 352046 500810 352102
rect 500878 352046 500934 352102
rect 501002 352046 501058 352102
rect 501126 352046 501182 352102
rect 500754 351922 500810 351978
rect 500878 351922 500934 351978
rect 501002 351922 501058 351978
rect 501126 351922 501182 351978
rect 502348 368702 502404 368758
rect 527754 364294 527810 364350
rect 527878 364294 527934 364350
rect 528002 364294 528058 364350
rect 528126 364294 528182 364350
rect 527754 364170 527810 364226
rect 527878 364170 527934 364226
rect 528002 364170 528058 364226
rect 528126 364170 528182 364226
rect 527754 364046 527810 364102
rect 527878 364046 527934 364102
rect 528002 364046 528058 364102
rect 528126 364046 528182 364102
rect 527754 363922 527810 363978
rect 527878 363922 527934 363978
rect 528002 363922 528058 363978
rect 528126 363922 528182 363978
rect 527754 346294 527810 346350
rect 527878 346294 527934 346350
rect 528002 346294 528058 346350
rect 528126 346294 528182 346350
rect 527754 346170 527810 346226
rect 527878 346170 527934 346226
rect 528002 346170 528058 346226
rect 528126 346170 528182 346226
rect 527754 346046 527810 346102
rect 527878 346046 527934 346102
rect 528002 346046 528058 346102
rect 528126 346046 528182 346102
rect 527754 345922 527810 345978
rect 527878 345922 527934 345978
rect 528002 345922 528058 345978
rect 528126 345922 528182 345978
rect 519484 345662 519540 345718
rect 516124 345482 516180 345538
rect 509404 345302 509460 345358
rect 512764 345122 512820 345178
rect 499878 334294 499934 334350
rect 500002 334294 500058 334350
rect 499878 334170 499934 334226
rect 500002 334170 500058 334226
rect 499878 334046 499934 334102
rect 500002 334046 500058 334102
rect 499878 333922 499934 333978
rect 500002 333922 500058 333978
rect 484518 328294 484574 328350
rect 484642 328294 484698 328350
rect 484518 328170 484574 328226
rect 484642 328170 484698 328226
rect 484518 328046 484574 328102
rect 484642 328046 484698 328102
rect 484518 327922 484574 327978
rect 484642 327922 484698 327978
rect 515238 328294 515294 328350
rect 515362 328294 515418 328350
rect 515238 328170 515294 328226
rect 515362 328170 515418 328226
rect 515238 328046 515294 328102
rect 515362 328046 515418 328102
rect 515238 327922 515294 327978
rect 515362 327922 515418 327978
rect 527754 328294 527810 328350
rect 527878 328294 527934 328350
rect 528002 328294 528058 328350
rect 528126 328294 528182 328350
rect 527754 328170 527810 328226
rect 527878 328170 527934 328226
rect 528002 328170 528058 328226
rect 528126 328170 528182 328226
rect 527754 328046 527810 328102
rect 527878 328046 527934 328102
rect 528002 328046 528058 328102
rect 528126 328046 528182 328102
rect 527754 327922 527810 327978
rect 527878 327922 527934 327978
rect 528002 327922 528058 327978
rect 528126 327922 528182 327978
rect 499878 316294 499934 316350
rect 500002 316294 500058 316350
rect 499878 316170 499934 316226
rect 500002 316170 500058 316226
rect 499878 316046 499934 316102
rect 500002 316046 500058 316102
rect 499878 315922 499934 315978
rect 500002 315922 500058 315978
rect 484518 310294 484574 310350
rect 484642 310294 484698 310350
rect 484518 310170 484574 310226
rect 484642 310170 484698 310226
rect 484518 310046 484574 310102
rect 484642 310046 484698 310102
rect 484518 309922 484574 309978
rect 484642 309922 484698 309978
rect 515238 310294 515294 310350
rect 515362 310294 515418 310350
rect 515238 310170 515294 310226
rect 515362 310170 515418 310226
rect 515238 310046 515294 310102
rect 515362 310046 515418 310102
rect 515238 309922 515294 309978
rect 515362 309922 515418 309978
rect 527754 310294 527810 310350
rect 527878 310294 527934 310350
rect 528002 310294 528058 310350
rect 528126 310294 528182 310350
rect 527754 310170 527810 310226
rect 527878 310170 527934 310226
rect 528002 310170 528058 310226
rect 528126 310170 528182 310226
rect 527754 310046 527810 310102
rect 527878 310046 527934 310102
rect 528002 310046 528058 310102
rect 528126 310046 528182 310102
rect 527754 309922 527810 309978
rect 527878 309922 527934 309978
rect 528002 309922 528058 309978
rect 528126 309922 528182 309978
rect 480172 298862 480228 298918
rect 480060 293822 480116 293878
rect 479836 283742 479892 283798
rect 497034 292294 497090 292350
rect 497158 292294 497214 292350
rect 497282 292294 497338 292350
rect 497406 292294 497462 292350
rect 497034 292170 497090 292226
rect 497158 292170 497214 292226
rect 497282 292170 497338 292226
rect 497406 292170 497462 292226
rect 497034 292046 497090 292102
rect 497158 292046 497214 292102
rect 497282 292046 497338 292102
rect 497406 292046 497462 292102
rect 497034 291922 497090 291978
rect 497158 291922 497214 291978
rect 497282 291922 497338 291978
rect 497406 291922 497462 291978
rect 497034 274294 497090 274350
rect 497158 274294 497214 274350
rect 497282 274294 497338 274350
rect 497406 274294 497462 274350
rect 497034 274170 497090 274226
rect 497158 274170 497214 274226
rect 497282 274170 497338 274226
rect 497406 274170 497462 274226
rect 497034 274046 497090 274102
rect 497158 274046 497214 274102
rect 497282 274046 497338 274102
rect 497406 274046 497462 274102
rect 497034 273922 497090 273978
rect 497158 273922 497214 273978
rect 497282 273922 497338 273978
rect 497406 273922 497462 273978
rect 470034 262294 470090 262350
rect 470158 262294 470214 262350
rect 470282 262294 470338 262350
rect 470406 262294 470462 262350
rect 470034 262170 470090 262226
rect 470158 262170 470214 262226
rect 470282 262170 470338 262226
rect 470406 262170 470462 262226
rect 470034 262046 470090 262102
rect 470158 262046 470214 262102
rect 470282 262046 470338 262102
rect 470406 262046 470462 262102
rect 470034 261922 470090 261978
rect 470158 261922 470214 261978
rect 470282 261922 470338 261978
rect 470406 261922 470462 261978
rect 497034 256294 497090 256350
rect 497158 256294 497214 256350
rect 497282 256294 497338 256350
rect 497406 256294 497462 256350
rect 497034 256170 497090 256226
rect 497158 256170 497214 256226
rect 497282 256170 497338 256226
rect 497406 256170 497462 256226
rect 497034 256046 497090 256102
rect 497158 256046 497214 256102
rect 497282 256046 497338 256102
rect 497406 256046 497462 256102
rect 472732 255967 472788 256023
rect 472856 255967 472912 256023
rect 472980 255967 473036 256023
rect 473104 255967 473160 256023
rect 472732 255843 472788 255899
rect 472856 255843 472912 255899
rect 472980 255843 473036 255899
rect 473104 255843 473160 255899
rect 497034 255922 497090 255978
rect 497158 255922 497214 255978
rect 497282 255922 497338 255978
rect 497406 255922 497462 255978
rect 470034 244294 470090 244350
rect 470158 244294 470214 244350
rect 470282 244294 470338 244350
rect 470406 244294 470462 244350
rect 470034 244170 470090 244226
rect 470158 244170 470214 244226
rect 470282 244170 470338 244226
rect 470406 244170 470462 244226
rect 470034 244046 470090 244102
rect 470158 244046 470214 244102
rect 470282 244046 470338 244102
rect 470406 244046 470462 244102
rect 470034 243922 470090 243978
rect 470158 243922 470214 243978
rect 470282 243922 470338 243978
rect 470406 243922 470462 243978
rect 471932 244294 471988 244350
rect 472056 244294 472112 244350
rect 472180 244294 472236 244350
rect 472304 244294 472360 244350
rect 471932 244170 471988 244226
rect 472056 244170 472112 244226
rect 472180 244170 472236 244226
rect 472304 244170 472360 244226
rect 471932 244046 471988 244102
rect 472056 244046 472112 244102
rect 472180 244046 472236 244102
rect 472304 244046 472360 244102
rect 471932 243922 471988 243978
rect 472056 243922 472112 243978
rect 472180 243922 472236 243978
rect 472304 243922 472360 243978
rect 472732 238294 472788 238350
rect 472856 238294 472912 238350
rect 472980 238294 473036 238350
rect 473104 238294 473160 238350
rect 472732 238170 472788 238226
rect 472856 238170 472912 238226
rect 472980 238170 473036 238226
rect 473104 238170 473160 238226
rect 472732 238046 472788 238102
rect 472856 238046 472912 238102
rect 472980 238046 473036 238102
rect 473104 238046 473160 238102
rect 472732 237922 472788 237978
rect 472856 237922 472912 237978
rect 472980 237922 473036 237978
rect 473104 237922 473160 237978
rect 497034 238294 497090 238350
rect 497158 238294 497214 238350
rect 497282 238294 497338 238350
rect 497406 238294 497462 238350
rect 497034 238170 497090 238226
rect 497158 238170 497214 238226
rect 497282 238170 497338 238226
rect 497406 238170 497462 238226
rect 497034 238046 497090 238102
rect 497158 238046 497214 238102
rect 497282 238046 497338 238102
rect 497406 238046 497462 238102
rect 497034 237922 497090 237978
rect 497158 237922 497214 237978
rect 497282 237922 497338 237978
rect 497406 237922 497462 237978
rect 470034 226294 470090 226350
rect 470158 226294 470214 226350
rect 470282 226294 470338 226350
rect 470406 226294 470462 226350
rect 470034 226170 470090 226226
rect 470158 226170 470214 226226
rect 470282 226170 470338 226226
rect 470406 226170 470462 226226
rect 470034 226046 470090 226102
rect 470158 226046 470214 226102
rect 470282 226046 470338 226102
rect 470406 226046 470462 226102
rect 470034 225922 470090 225978
rect 470158 225922 470214 225978
rect 470282 225922 470338 225978
rect 470406 225922 470462 225978
rect 471932 226294 471988 226350
rect 472056 226294 472112 226350
rect 472180 226294 472236 226350
rect 472304 226294 472360 226350
rect 471932 226170 471988 226226
rect 472056 226170 472112 226226
rect 472180 226170 472236 226226
rect 472304 226170 472360 226226
rect 471932 226046 471988 226102
rect 472056 226046 472112 226102
rect 472180 226046 472236 226102
rect 472304 226046 472360 226102
rect 471932 225922 471988 225978
rect 472056 225922 472112 225978
rect 472180 225922 472236 225978
rect 472304 225922 472360 225978
rect 472732 220294 472788 220350
rect 472856 220294 472912 220350
rect 472980 220294 473036 220350
rect 473104 220294 473160 220350
rect 472732 220170 472788 220226
rect 472856 220170 472912 220226
rect 472980 220170 473036 220226
rect 473104 220170 473160 220226
rect 472732 220046 472788 220102
rect 472856 220046 472912 220102
rect 472980 220046 473036 220102
rect 473104 220046 473160 220102
rect 472732 219922 472788 219978
rect 472856 219922 472912 219978
rect 472980 219922 473036 219978
rect 473104 219922 473160 219978
rect 497034 220294 497090 220350
rect 497158 220294 497214 220350
rect 497282 220294 497338 220350
rect 497406 220294 497462 220350
rect 497034 220170 497090 220226
rect 497158 220170 497214 220226
rect 497282 220170 497338 220226
rect 497406 220170 497462 220226
rect 497034 220046 497090 220102
rect 497158 220046 497214 220102
rect 497282 220046 497338 220102
rect 497406 220046 497462 220102
rect 497034 219922 497090 219978
rect 497158 219922 497214 219978
rect 497282 219922 497338 219978
rect 497406 219922 497462 219978
rect 470034 208294 470090 208350
rect 470158 208294 470214 208350
rect 470282 208294 470338 208350
rect 470406 208294 470462 208350
rect 470034 208170 470090 208226
rect 470158 208170 470214 208226
rect 470282 208170 470338 208226
rect 470406 208170 470462 208226
rect 470034 208046 470090 208102
rect 470158 208046 470214 208102
rect 470282 208046 470338 208102
rect 470406 208046 470462 208102
rect 470034 207922 470090 207978
rect 470158 207922 470214 207978
rect 470282 207922 470338 207978
rect 470406 207922 470462 207978
rect 471932 208294 471988 208350
rect 472056 208294 472112 208350
rect 472180 208294 472236 208350
rect 472304 208294 472360 208350
rect 471932 208170 471988 208226
rect 472056 208170 472112 208226
rect 472180 208170 472236 208226
rect 472304 208170 472360 208226
rect 471932 208046 471988 208102
rect 472056 208046 472112 208102
rect 472180 208046 472236 208102
rect 472304 208046 472360 208102
rect 471932 207922 471988 207978
rect 472056 207922 472112 207978
rect 472180 207922 472236 207978
rect 472304 207922 472360 207978
rect 472732 202294 472788 202350
rect 472856 202294 472912 202350
rect 472980 202294 473036 202350
rect 473104 202294 473160 202350
rect 472732 202170 472788 202226
rect 472856 202170 472912 202226
rect 472980 202170 473036 202226
rect 473104 202170 473160 202226
rect 472732 202046 472788 202102
rect 472856 202046 472912 202102
rect 472980 202046 473036 202102
rect 473104 202046 473160 202102
rect 472732 201922 472788 201978
rect 472856 201922 472912 201978
rect 472980 201922 473036 201978
rect 473104 201922 473160 201978
rect 497034 202294 497090 202350
rect 497158 202294 497214 202350
rect 497282 202294 497338 202350
rect 497406 202294 497462 202350
rect 497034 202170 497090 202226
rect 497158 202170 497214 202226
rect 497282 202170 497338 202226
rect 497406 202170 497462 202226
rect 497034 202046 497090 202102
rect 497158 202046 497214 202102
rect 497282 202046 497338 202102
rect 497406 202046 497462 202102
rect 497034 201922 497090 201978
rect 497158 201922 497214 201978
rect 497282 201922 497338 201978
rect 497406 201922 497462 201978
rect 470034 190294 470090 190350
rect 470158 190294 470214 190350
rect 470282 190294 470338 190350
rect 470406 190294 470462 190350
rect 470034 190170 470090 190226
rect 470158 190170 470214 190226
rect 470282 190170 470338 190226
rect 470406 190170 470462 190226
rect 470034 190046 470090 190102
rect 470158 190046 470214 190102
rect 470282 190046 470338 190102
rect 470406 190046 470462 190102
rect 470034 189922 470090 189978
rect 470158 189922 470214 189978
rect 470282 189922 470338 189978
rect 470406 189922 470462 189978
rect 471932 190294 471988 190350
rect 472056 190294 472112 190350
rect 472180 190294 472236 190350
rect 472304 190294 472360 190350
rect 471932 190170 471988 190226
rect 472056 190170 472112 190226
rect 472180 190170 472236 190226
rect 472304 190170 472360 190226
rect 471932 190046 471988 190102
rect 472056 190046 472112 190102
rect 472180 190046 472236 190102
rect 472304 190046 472360 190102
rect 471932 189922 471988 189978
rect 472056 189922 472112 189978
rect 472180 189922 472236 189978
rect 472304 189922 472360 189978
rect 472732 184294 472788 184350
rect 472856 184294 472912 184350
rect 472980 184294 473036 184350
rect 473104 184294 473160 184350
rect 472732 184170 472788 184226
rect 472856 184170 472912 184226
rect 472980 184170 473036 184226
rect 473104 184170 473160 184226
rect 472732 184046 472788 184102
rect 472856 184046 472912 184102
rect 472980 184046 473036 184102
rect 473104 184046 473160 184102
rect 472732 183922 472788 183978
rect 472856 183922 472912 183978
rect 472980 183922 473036 183978
rect 473104 183922 473160 183978
rect 497034 184294 497090 184350
rect 497158 184294 497214 184350
rect 497282 184294 497338 184350
rect 497406 184294 497462 184350
rect 497034 184170 497090 184226
rect 497158 184170 497214 184226
rect 497282 184170 497338 184226
rect 497406 184170 497462 184226
rect 497034 184046 497090 184102
rect 497158 184046 497214 184102
rect 497282 184046 497338 184102
rect 497406 184046 497462 184102
rect 497034 183922 497090 183978
rect 497158 183922 497214 183978
rect 497282 183922 497338 183978
rect 497406 183922 497462 183978
rect 470034 172294 470090 172350
rect 470158 172294 470214 172350
rect 470282 172294 470338 172350
rect 470406 172294 470462 172350
rect 470034 172170 470090 172226
rect 470158 172170 470214 172226
rect 470282 172170 470338 172226
rect 470406 172170 470462 172226
rect 470034 172046 470090 172102
rect 470158 172046 470214 172102
rect 470282 172046 470338 172102
rect 470406 172046 470462 172102
rect 470034 171922 470090 171978
rect 470158 171922 470214 171978
rect 470282 171922 470338 171978
rect 470406 171922 470462 171978
rect 471932 172294 471988 172350
rect 472056 172294 472112 172350
rect 472180 172294 472236 172350
rect 472304 172294 472360 172350
rect 471932 172170 471988 172226
rect 472056 172170 472112 172226
rect 472180 172170 472236 172226
rect 472304 172170 472360 172226
rect 471932 172046 471988 172102
rect 472056 172046 472112 172102
rect 472180 172046 472236 172102
rect 472304 172046 472360 172102
rect 471932 171922 471988 171978
rect 472056 171922 472112 171978
rect 472180 171922 472236 171978
rect 472304 171922 472360 171978
rect 472732 166294 472788 166350
rect 472856 166294 472912 166350
rect 472980 166294 473036 166350
rect 473104 166294 473160 166350
rect 472732 166170 472788 166226
rect 472856 166170 472912 166226
rect 472980 166170 473036 166226
rect 473104 166170 473160 166226
rect 472732 166046 472788 166102
rect 472856 166046 472912 166102
rect 472980 166046 473036 166102
rect 473104 166046 473160 166102
rect 472732 165922 472788 165978
rect 472856 165922 472912 165978
rect 472980 165922 473036 165978
rect 473104 165922 473160 165978
rect 497034 166294 497090 166350
rect 497158 166294 497214 166350
rect 497282 166294 497338 166350
rect 497406 166294 497462 166350
rect 497034 166170 497090 166226
rect 497158 166170 497214 166226
rect 497282 166170 497338 166226
rect 497406 166170 497462 166226
rect 497034 166046 497090 166102
rect 497158 166046 497214 166102
rect 497282 166046 497338 166102
rect 497406 166046 497462 166102
rect 497034 165922 497090 165978
rect 497158 165922 497214 165978
rect 497282 165922 497338 165978
rect 497406 165922 497462 165978
rect 470034 154294 470090 154350
rect 470158 154294 470214 154350
rect 470282 154294 470338 154350
rect 470406 154294 470462 154350
rect 470034 154170 470090 154226
rect 470158 154170 470214 154226
rect 470282 154170 470338 154226
rect 470406 154170 470462 154226
rect 470034 154046 470090 154102
rect 470158 154046 470214 154102
rect 470282 154046 470338 154102
rect 470406 154046 470462 154102
rect 470034 153922 470090 153978
rect 470158 153922 470214 153978
rect 470282 153922 470338 153978
rect 470406 153922 470462 153978
rect 474572 142442 474628 142498
rect 497034 148294 497090 148350
rect 497158 148294 497214 148350
rect 497282 148294 497338 148350
rect 497406 148294 497462 148350
rect 497034 148170 497090 148226
rect 497158 148170 497214 148226
rect 497282 148170 497338 148226
rect 497406 148170 497462 148226
rect 497034 148046 497090 148102
rect 497158 148046 497214 148102
rect 497282 148046 497338 148102
rect 497406 148046 497462 148102
rect 497034 147922 497090 147978
rect 497158 147922 497214 147978
rect 497282 147922 497338 147978
rect 497406 147922 497462 147978
rect 471996 142262 472052 142318
rect 484428 141902 484484 141958
rect 470034 136294 470090 136350
rect 470158 136294 470214 136350
rect 470282 136294 470338 136350
rect 470406 136294 470462 136350
rect 470034 136170 470090 136226
rect 470158 136170 470214 136226
rect 470282 136170 470338 136226
rect 470406 136170 470462 136226
rect 470034 136046 470090 136102
rect 470158 136046 470214 136102
rect 470282 136046 470338 136102
rect 470406 136046 470462 136102
rect 470034 135922 470090 135978
rect 470158 135922 470214 135978
rect 470282 135922 470338 135978
rect 470406 135922 470462 135978
rect 470034 118294 470090 118350
rect 470158 118294 470214 118350
rect 470282 118294 470338 118350
rect 470406 118294 470462 118350
rect 470034 118170 470090 118226
rect 470158 118170 470214 118226
rect 470282 118170 470338 118226
rect 470406 118170 470462 118226
rect 470034 118046 470090 118102
rect 470158 118046 470214 118102
rect 470282 118046 470338 118102
rect 470406 118046 470462 118102
rect 470034 117922 470090 117978
rect 470158 117922 470214 117978
rect 470282 117922 470338 117978
rect 470406 117922 470462 117978
rect 470034 100294 470090 100350
rect 470158 100294 470214 100350
rect 470282 100294 470338 100350
rect 470406 100294 470462 100350
rect 470034 100170 470090 100226
rect 470158 100170 470214 100226
rect 470282 100170 470338 100226
rect 470406 100170 470462 100226
rect 470034 100046 470090 100102
rect 470158 100046 470214 100102
rect 470282 100046 470338 100102
rect 470406 100046 470462 100102
rect 470034 99922 470090 99978
rect 470158 99922 470214 99978
rect 470282 99922 470338 99978
rect 470406 99922 470462 99978
rect 470034 82294 470090 82350
rect 470158 82294 470214 82350
rect 470282 82294 470338 82350
rect 470406 82294 470462 82350
rect 470034 82170 470090 82226
rect 470158 82170 470214 82226
rect 470282 82170 470338 82226
rect 470406 82170 470462 82226
rect 470034 82046 470090 82102
rect 470158 82046 470214 82102
rect 470282 82046 470338 82102
rect 470406 82046 470462 82102
rect 470034 81922 470090 81978
rect 470158 81922 470214 81978
rect 470282 81922 470338 81978
rect 470406 81922 470462 81978
rect 470034 64294 470090 64350
rect 470158 64294 470214 64350
rect 470282 64294 470338 64350
rect 470406 64294 470462 64350
rect 470034 64170 470090 64226
rect 470158 64170 470214 64226
rect 470282 64170 470338 64226
rect 470406 64170 470462 64226
rect 470034 64046 470090 64102
rect 470158 64046 470214 64102
rect 470282 64046 470338 64102
rect 470406 64046 470462 64102
rect 470034 63922 470090 63978
rect 470158 63922 470214 63978
rect 470282 63922 470338 63978
rect 470406 63922 470462 63978
rect 470034 46294 470090 46350
rect 470158 46294 470214 46350
rect 470282 46294 470338 46350
rect 470406 46294 470462 46350
rect 470034 46170 470090 46226
rect 470158 46170 470214 46226
rect 470282 46170 470338 46226
rect 470406 46170 470462 46226
rect 470034 46046 470090 46102
rect 470158 46046 470214 46102
rect 470282 46046 470338 46102
rect 470406 46046 470462 46102
rect 470034 45922 470090 45978
rect 470158 45922 470214 45978
rect 470282 45922 470338 45978
rect 470406 45922 470462 45978
rect 470034 28294 470090 28350
rect 470158 28294 470214 28350
rect 470282 28294 470338 28350
rect 470406 28294 470462 28350
rect 470034 28170 470090 28226
rect 470158 28170 470214 28226
rect 470282 28170 470338 28226
rect 470406 28170 470462 28226
rect 470034 28046 470090 28102
rect 470158 28046 470214 28102
rect 470282 28046 470338 28102
rect 470406 28046 470462 28102
rect 470034 27922 470090 27978
rect 470158 27922 470214 27978
rect 470282 27922 470338 27978
rect 470406 27922 470462 27978
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 500754 298294 500810 298350
rect 500878 298294 500934 298350
rect 501002 298294 501058 298350
rect 501126 298294 501182 298350
rect 500754 298170 500810 298226
rect 500878 298170 500934 298226
rect 501002 298170 501058 298226
rect 501126 298170 501182 298226
rect 500754 298046 500810 298102
rect 500878 298046 500934 298102
rect 501002 298046 501058 298102
rect 501126 298046 501182 298102
rect 500754 297922 500810 297978
rect 500878 297922 500934 297978
rect 501002 297922 501058 297978
rect 501126 297922 501182 297978
rect 500754 280294 500810 280350
rect 500878 280294 500934 280350
rect 501002 280294 501058 280350
rect 501126 280294 501182 280350
rect 500754 280170 500810 280226
rect 500878 280170 500934 280226
rect 501002 280170 501058 280226
rect 501126 280170 501182 280226
rect 500754 280046 500810 280102
rect 500878 280046 500934 280102
rect 501002 280046 501058 280102
rect 501126 280046 501182 280102
rect 500754 279922 500810 279978
rect 500878 279922 500934 279978
rect 501002 279922 501058 279978
rect 501126 279922 501182 279978
rect 500754 262294 500810 262350
rect 500878 262294 500934 262350
rect 501002 262294 501058 262350
rect 501126 262294 501182 262350
rect 500754 262170 500810 262226
rect 500878 262170 500934 262226
rect 501002 262170 501058 262226
rect 501126 262170 501182 262226
rect 500754 262046 500810 262102
rect 500878 262046 500934 262102
rect 501002 262046 501058 262102
rect 501126 262046 501182 262102
rect 500754 261922 500810 261978
rect 500878 261922 500934 261978
rect 501002 261922 501058 261978
rect 501126 261922 501182 261978
rect 500754 244294 500810 244350
rect 500878 244294 500934 244350
rect 501002 244294 501058 244350
rect 501126 244294 501182 244350
rect 500754 244170 500810 244226
rect 500878 244170 500934 244226
rect 501002 244170 501058 244226
rect 501126 244170 501182 244226
rect 500754 244046 500810 244102
rect 500878 244046 500934 244102
rect 501002 244046 501058 244102
rect 501126 244046 501182 244102
rect 500754 243922 500810 243978
rect 500878 243922 500934 243978
rect 501002 243922 501058 243978
rect 501126 243922 501182 243978
rect 500754 226294 500810 226350
rect 500878 226294 500934 226350
rect 501002 226294 501058 226350
rect 501126 226294 501182 226350
rect 500754 226170 500810 226226
rect 500878 226170 500934 226226
rect 501002 226170 501058 226226
rect 501126 226170 501182 226226
rect 500754 226046 500810 226102
rect 500878 226046 500934 226102
rect 501002 226046 501058 226102
rect 501126 226046 501182 226102
rect 500754 225922 500810 225978
rect 500878 225922 500934 225978
rect 501002 225922 501058 225978
rect 501126 225922 501182 225978
rect 500754 208294 500810 208350
rect 500878 208294 500934 208350
rect 501002 208294 501058 208350
rect 501126 208294 501182 208350
rect 500754 208170 500810 208226
rect 500878 208170 500934 208226
rect 501002 208170 501058 208226
rect 501126 208170 501182 208226
rect 500754 208046 500810 208102
rect 500878 208046 500934 208102
rect 501002 208046 501058 208102
rect 501126 208046 501182 208102
rect 500754 207922 500810 207978
rect 500878 207922 500934 207978
rect 501002 207922 501058 207978
rect 501126 207922 501182 207978
rect 500754 190294 500810 190350
rect 500878 190294 500934 190350
rect 501002 190294 501058 190350
rect 501126 190294 501182 190350
rect 500754 190170 500810 190226
rect 500878 190170 500934 190226
rect 501002 190170 501058 190226
rect 501126 190170 501182 190226
rect 500754 190046 500810 190102
rect 500878 190046 500934 190102
rect 501002 190046 501058 190102
rect 501126 190046 501182 190102
rect 500754 189922 500810 189978
rect 500878 189922 500934 189978
rect 501002 189922 501058 189978
rect 501126 189922 501182 189978
rect 500754 172294 500810 172350
rect 500878 172294 500934 172350
rect 501002 172294 501058 172350
rect 501126 172294 501182 172350
rect 500754 172170 500810 172226
rect 500878 172170 500934 172226
rect 501002 172170 501058 172226
rect 501126 172170 501182 172226
rect 500754 172046 500810 172102
rect 500878 172046 500934 172102
rect 501002 172046 501058 172102
rect 501126 172046 501182 172102
rect 500754 171922 500810 171978
rect 500878 171922 500934 171978
rect 501002 171922 501058 171978
rect 501126 171922 501182 171978
rect 500754 154294 500810 154350
rect 500878 154294 500934 154350
rect 501002 154294 501058 154350
rect 501126 154294 501182 154350
rect 500754 154170 500810 154226
rect 500878 154170 500934 154226
rect 501002 154170 501058 154226
rect 501126 154170 501182 154226
rect 500754 154046 500810 154102
rect 500878 154046 500934 154102
rect 501002 154046 501058 154102
rect 501126 154046 501182 154102
rect 500754 153922 500810 153978
rect 500878 153922 500934 153978
rect 501002 153922 501058 153978
rect 501126 153922 501182 153978
rect 498988 142622 499044 142678
rect 497034 130294 497090 130350
rect 497158 130294 497214 130350
rect 497282 130294 497338 130350
rect 497406 130294 497462 130350
rect 497034 130170 497090 130226
rect 497158 130170 497214 130226
rect 497282 130170 497338 130226
rect 497406 130170 497462 130226
rect 497034 130046 497090 130102
rect 497158 130046 497214 130102
rect 497282 130046 497338 130102
rect 497406 130046 497462 130102
rect 497034 129922 497090 129978
rect 497158 129922 497214 129978
rect 497282 129922 497338 129978
rect 497406 129922 497462 129978
rect 497034 112294 497090 112350
rect 497158 112294 497214 112350
rect 497282 112294 497338 112350
rect 497406 112294 497462 112350
rect 497034 112170 497090 112226
rect 497158 112170 497214 112226
rect 497282 112170 497338 112226
rect 497406 112170 497462 112226
rect 497034 112046 497090 112102
rect 497158 112046 497214 112102
rect 497282 112046 497338 112102
rect 497406 112046 497462 112102
rect 497034 111922 497090 111978
rect 497158 111922 497214 111978
rect 497282 111922 497338 111978
rect 497406 111922 497462 111978
rect 497034 94294 497090 94350
rect 497158 94294 497214 94350
rect 497282 94294 497338 94350
rect 497406 94294 497462 94350
rect 497034 94170 497090 94226
rect 497158 94170 497214 94226
rect 497282 94170 497338 94226
rect 497406 94170 497462 94226
rect 497034 94046 497090 94102
rect 497158 94046 497214 94102
rect 497282 94046 497338 94102
rect 497406 94046 497462 94102
rect 497034 93922 497090 93978
rect 497158 93922 497214 93978
rect 497282 93922 497338 93978
rect 497406 93922 497462 93978
rect 497034 76294 497090 76350
rect 497158 76294 497214 76350
rect 497282 76294 497338 76350
rect 497406 76294 497462 76350
rect 497034 76170 497090 76226
rect 497158 76170 497214 76226
rect 497282 76170 497338 76226
rect 497406 76170 497462 76226
rect 497034 76046 497090 76102
rect 497158 76046 497214 76102
rect 497282 76046 497338 76102
rect 497406 76046 497462 76102
rect 497034 75922 497090 75978
rect 497158 75922 497214 75978
rect 497282 75922 497338 75978
rect 497406 75922 497462 75978
rect 497034 58294 497090 58350
rect 497158 58294 497214 58350
rect 497282 58294 497338 58350
rect 497406 58294 497462 58350
rect 497034 58170 497090 58226
rect 497158 58170 497214 58226
rect 497282 58170 497338 58226
rect 497406 58170 497462 58226
rect 497034 58046 497090 58102
rect 497158 58046 497214 58102
rect 497282 58046 497338 58102
rect 497406 58046 497462 58102
rect 497034 57922 497090 57978
rect 497158 57922 497214 57978
rect 497282 57922 497338 57978
rect 497406 57922 497462 57978
rect 497034 40294 497090 40350
rect 497158 40294 497214 40350
rect 497282 40294 497338 40350
rect 497406 40294 497462 40350
rect 497034 40170 497090 40226
rect 497158 40170 497214 40226
rect 497282 40170 497338 40226
rect 497406 40170 497462 40226
rect 497034 40046 497090 40102
rect 497158 40046 497214 40102
rect 497282 40046 497338 40102
rect 497406 40046 497462 40102
rect 497034 39922 497090 39978
rect 497158 39922 497214 39978
rect 497282 39922 497338 39978
rect 497406 39922 497462 39978
rect 497034 22294 497090 22350
rect 497158 22294 497214 22350
rect 497282 22294 497338 22350
rect 497406 22294 497462 22350
rect 497034 22170 497090 22226
rect 497158 22170 497214 22226
rect 497282 22170 497338 22226
rect 497406 22170 497462 22226
rect 497034 22046 497090 22102
rect 497158 22046 497214 22102
rect 497282 22046 497338 22102
rect 497406 22046 497462 22102
rect 497034 21922 497090 21978
rect 497158 21922 497214 21978
rect 497282 21922 497338 21978
rect 497406 21922 497462 21978
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 527754 292294 527810 292350
rect 527878 292294 527934 292350
rect 528002 292294 528058 292350
rect 528126 292294 528182 292350
rect 527754 292170 527810 292226
rect 527878 292170 527934 292226
rect 528002 292170 528058 292226
rect 528126 292170 528182 292226
rect 527754 292046 527810 292102
rect 527878 292046 527934 292102
rect 528002 292046 528058 292102
rect 528126 292046 528182 292102
rect 527754 291922 527810 291978
rect 527878 291922 527934 291978
rect 528002 291922 528058 291978
rect 528126 291922 528182 291978
rect 527754 274294 527810 274350
rect 527878 274294 527934 274350
rect 528002 274294 528058 274350
rect 528126 274294 528182 274350
rect 527754 274170 527810 274226
rect 527878 274170 527934 274226
rect 528002 274170 528058 274226
rect 528126 274170 528182 274226
rect 527754 274046 527810 274102
rect 527878 274046 527934 274102
rect 528002 274046 528058 274102
rect 528126 274046 528182 274102
rect 527754 273922 527810 273978
rect 527878 273922 527934 273978
rect 528002 273922 528058 273978
rect 528126 273922 528182 273978
rect 527754 256294 527810 256350
rect 527878 256294 527934 256350
rect 528002 256294 528058 256350
rect 528126 256294 528182 256350
rect 527754 256170 527810 256226
rect 527878 256170 527934 256226
rect 528002 256170 528058 256226
rect 528126 256170 528182 256226
rect 527754 256046 527810 256102
rect 527878 256046 527934 256102
rect 528002 256046 528058 256102
rect 528126 256046 528182 256102
rect 527754 255922 527810 255978
rect 527878 255922 527934 255978
rect 528002 255922 528058 255978
rect 528126 255922 528182 255978
rect 527754 238294 527810 238350
rect 527878 238294 527934 238350
rect 528002 238294 528058 238350
rect 528126 238294 528182 238350
rect 527754 238170 527810 238226
rect 527878 238170 527934 238226
rect 528002 238170 528058 238226
rect 528126 238170 528182 238226
rect 527754 238046 527810 238102
rect 527878 238046 527934 238102
rect 528002 238046 528058 238102
rect 528126 238046 528182 238102
rect 527754 237922 527810 237978
rect 527878 237922 527934 237978
rect 528002 237922 528058 237978
rect 528126 237922 528182 237978
rect 527754 220294 527810 220350
rect 527878 220294 527934 220350
rect 528002 220294 528058 220350
rect 528126 220294 528182 220350
rect 527754 220170 527810 220226
rect 527878 220170 527934 220226
rect 528002 220170 528058 220226
rect 528126 220170 528182 220226
rect 527754 220046 527810 220102
rect 527878 220046 527934 220102
rect 528002 220046 528058 220102
rect 528126 220046 528182 220102
rect 527754 219922 527810 219978
rect 527878 219922 527934 219978
rect 528002 219922 528058 219978
rect 528126 219922 528182 219978
rect 527754 202294 527810 202350
rect 527878 202294 527934 202350
rect 528002 202294 528058 202350
rect 528126 202294 528182 202350
rect 527754 202170 527810 202226
rect 527878 202170 527934 202226
rect 528002 202170 528058 202226
rect 528126 202170 528182 202226
rect 527754 202046 527810 202102
rect 527878 202046 527934 202102
rect 528002 202046 528058 202102
rect 528126 202046 528182 202102
rect 527754 201922 527810 201978
rect 527878 201922 527934 201978
rect 528002 201922 528058 201978
rect 528126 201922 528182 201978
rect 527754 184294 527810 184350
rect 527878 184294 527934 184350
rect 528002 184294 528058 184350
rect 528126 184294 528182 184350
rect 527754 184170 527810 184226
rect 527878 184170 527934 184226
rect 528002 184170 528058 184226
rect 528126 184170 528182 184226
rect 527754 184046 527810 184102
rect 527878 184046 527934 184102
rect 528002 184046 528058 184102
rect 528126 184046 528182 184102
rect 527754 183922 527810 183978
rect 527878 183922 527934 183978
rect 528002 183922 528058 183978
rect 528126 183922 528182 183978
rect 527754 166294 527810 166350
rect 527878 166294 527934 166350
rect 528002 166294 528058 166350
rect 528126 166294 528182 166350
rect 527754 166170 527810 166226
rect 527878 166170 527934 166226
rect 528002 166170 528058 166226
rect 528126 166170 528182 166226
rect 527754 166046 527810 166102
rect 527878 166046 527934 166102
rect 528002 166046 528058 166102
rect 528126 166046 528182 166102
rect 527754 165922 527810 165978
rect 527878 165922 527934 165978
rect 528002 165922 528058 165978
rect 528126 165922 528182 165978
rect 527754 148294 527810 148350
rect 527878 148294 527934 148350
rect 528002 148294 528058 148350
rect 528126 148294 528182 148350
rect 527754 148170 527810 148226
rect 527878 148170 527934 148226
rect 528002 148170 528058 148226
rect 528126 148170 528182 148226
rect 527754 148046 527810 148102
rect 527878 148046 527934 148102
rect 528002 148046 528058 148102
rect 528126 148046 528182 148102
rect 527754 147922 527810 147978
rect 527878 147922 527934 147978
rect 528002 147922 528058 147978
rect 528126 147922 528182 147978
rect 505596 141002 505652 141058
rect 500754 136294 500810 136350
rect 500878 136294 500934 136350
rect 501002 136294 501058 136350
rect 501126 136294 501182 136350
rect 500754 136170 500810 136226
rect 500878 136170 500934 136226
rect 501002 136170 501058 136226
rect 501126 136170 501182 136226
rect 500754 136046 500810 136102
rect 500878 136046 500934 136102
rect 501002 136046 501058 136102
rect 501126 136046 501182 136102
rect 500754 135922 500810 135978
rect 500878 135922 500934 135978
rect 501002 135922 501058 135978
rect 501126 135922 501182 135978
rect 500754 118294 500810 118350
rect 500878 118294 500934 118350
rect 501002 118294 501058 118350
rect 501126 118294 501182 118350
rect 500754 118170 500810 118226
rect 500878 118170 500934 118226
rect 501002 118170 501058 118226
rect 501126 118170 501182 118226
rect 500754 118046 500810 118102
rect 500878 118046 500934 118102
rect 501002 118046 501058 118102
rect 501126 118046 501182 118102
rect 500754 117922 500810 117978
rect 500878 117922 500934 117978
rect 501002 117922 501058 117978
rect 501126 117922 501182 117978
rect 500754 100294 500810 100350
rect 500878 100294 500934 100350
rect 501002 100294 501058 100350
rect 501126 100294 501182 100350
rect 500754 100170 500810 100226
rect 500878 100170 500934 100226
rect 501002 100170 501058 100226
rect 501126 100170 501182 100226
rect 500754 100046 500810 100102
rect 500878 100046 500934 100102
rect 501002 100046 501058 100102
rect 501126 100046 501182 100102
rect 500754 99922 500810 99978
rect 500878 99922 500934 99978
rect 501002 99922 501058 99978
rect 501126 99922 501182 99978
rect 500754 82294 500810 82350
rect 500878 82294 500934 82350
rect 501002 82294 501058 82350
rect 501126 82294 501182 82350
rect 500754 82170 500810 82226
rect 500878 82170 500934 82226
rect 501002 82170 501058 82226
rect 501126 82170 501182 82226
rect 500754 82046 500810 82102
rect 500878 82046 500934 82102
rect 501002 82046 501058 82102
rect 501126 82046 501182 82102
rect 500754 81922 500810 81978
rect 500878 81922 500934 81978
rect 501002 81922 501058 81978
rect 501126 81922 501182 81978
rect 500754 64294 500810 64350
rect 500878 64294 500934 64350
rect 501002 64294 501058 64350
rect 501126 64294 501182 64350
rect 500754 64170 500810 64226
rect 500878 64170 500934 64226
rect 501002 64170 501058 64226
rect 501126 64170 501182 64226
rect 500754 64046 500810 64102
rect 500878 64046 500934 64102
rect 501002 64046 501058 64102
rect 501126 64046 501182 64102
rect 500754 63922 500810 63978
rect 500878 63922 500934 63978
rect 501002 63922 501058 63978
rect 501126 63922 501182 63978
rect 500754 46294 500810 46350
rect 500878 46294 500934 46350
rect 501002 46294 501058 46350
rect 501126 46294 501182 46350
rect 500754 46170 500810 46226
rect 500878 46170 500934 46226
rect 501002 46170 501058 46226
rect 501126 46170 501182 46226
rect 500754 46046 500810 46102
rect 500878 46046 500934 46102
rect 501002 46046 501058 46102
rect 501126 46046 501182 46102
rect 500754 45922 500810 45978
rect 500878 45922 500934 45978
rect 501002 45922 501058 45978
rect 501126 45922 501182 45978
rect 500754 28294 500810 28350
rect 500878 28294 500934 28350
rect 501002 28294 501058 28350
rect 501126 28294 501182 28350
rect 500754 28170 500810 28226
rect 500878 28170 500934 28226
rect 501002 28170 501058 28226
rect 501126 28170 501182 28226
rect 500754 28046 500810 28102
rect 500878 28046 500934 28102
rect 501002 28046 501058 28102
rect 501126 28046 501182 28102
rect 500754 27922 500810 27978
rect 500878 27922 500934 27978
rect 501002 27922 501058 27978
rect 501126 27922 501182 27978
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 527754 130294 527810 130350
rect 527878 130294 527934 130350
rect 528002 130294 528058 130350
rect 528126 130294 528182 130350
rect 527754 130170 527810 130226
rect 527878 130170 527934 130226
rect 528002 130170 528058 130226
rect 528126 130170 528182 130226
rect 527754 130046 527810 130102
rect 527878 130046 527934 130102
rect 528002 130046 528058 130102
rect 528126 130046 528182 130102
rect 527754 129922 527810 129978
rect 527878 129922 527934 129978
rect 528002 129922 528058 129978
rect 528126 129922 528182 129978
rect 527754 112294 527810 112350
rect 527878 112294 527934 112350
rect 528002 112294 528058 112350
rect 528126 112294 528182 112350
rect 527754 112170 527810 112226
rect 527878 112170 527934 112226
rect 528002 112170 528058 112226
rect 528126 112170 528182 112226
rect 527754 112046 527810 112102
rect 527878 112046 527934 112102
rect 528002 112046 528058 112102
rect 528126 112046 528182 112102
rect 527754 111922 527810 111978
rect 527878 111922 527934 111978
rect 528002 111922 528058 111978
rect 528126 111922 528182 111978
rect 527754 94294 527810 94350
rect 527878 94294 527934 94350
rect 528002 94294 528058 94350
rect 528126 94294 528182 94350
rect 527754 94170 527810 94226
rect 527878 94170 527934 94226
rect 528002 94170 528058 94226
rect 528126 94170 528182 94226
rect 527754 94046 527810 94102
rect 527878 94046 527934 94102
rect 528002 94046 528058 94102
rect 528126 94046 528182 94102
rect 527754 93922 527810 93978
rect 527878 93922 527934 93978
rect 528002 93922 528058 93978
rect 528126 93922 528182 93978
rect 527754 76294 527810 76350
rect 527878 76294 527934 76350
rect 528002 76294 528058 76350
rect 528126 76294 528182 76350
rect 527754 76170 527810 76226
rect 527878 76170 527934 76226
rect 528002 76170 528058 76226
rect 528126 76170 528182 76226
rect 527754 76046 527810 76102
rect 527878 76046 527934 76102
rect 528002 76046 528058 76102
rect 528126 76046 528182 76102
rect 527754 75922 527810 75978
rect 527878 75922 527934 75978
rect 528002 75922 528058 75978
rect 528126 75922 528182 75978
rect 527754 58294 527810 58350
rect 527878 58294 527934 58350
rect 528002 58294 528058 58350
rect 528126 58294 528182 58350
rect 527754 58170 527810 58226
rect 527878 58170 527934 58226
rect 528002 58170 528058 58226
rect 528126 58170 528182 58226
rect 527754 58046 527810 58102
rect 527878 58046 527934 58102
rect 528002 58046 528058 58102
rect 528126 58046 528182 58102
rect 527754 57922 527810 57978
rect 527878 57922 527934 57978
rect 528002 57922 528058 57978
rect 528126 57922 528182 57978
rect 527754 40294 527810 40350
rect 527878 40294 527934 40350
rect 528002 40294 528058 40350
rect 528126 40294 528182 40350
rect 527754 40170 527810 40226
rect 527878 40170 527934 40226
rect 528002 40170 528058 40226
rect 528126 40170 528182 40226
rect 527754 40046 527810 40102
rect 527878 40046 527934 40102
rect 528002 40046 528058 40102
rect 528126 40046 528182 40102
rect 527754 39922 527810 39978
rect 527878 39922 527934 39978
rect 528002 39922 528058 39978
rect 528126 39922 528182 39978
rect 527754 22294 527810 22350
rect 527878 22294 527934 22350
rect 528002 22294 528058 22350
rect 528126 22294 528182 22350
rect 527754 22170 527810 22226
rect 527878 22170 527934 22226
rect 528002 22170 528058 22226
rect 528126 22170 528182 22226
rect 527754 22046 527810 22102
rect 527878 22046 527934 22102
rect 528002 22046 528058 22102
rect 528126 22046 528182 22102
rect 527754 21922 527810 21978
rect 527878 21922 527934 21978
rect 528002 21922 528058 21978
rect 528126 21922 528182 21978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 531474 442294 531530 442350
rect 531598 442294 531654 442350
rect 531722 442294 531778 442350
rect 531846 442294 531902 442350
rect 531474 442170 531530 442226
rect 531598 442170 531654 442226
rect 531722 442170 531778 442226
rect 531846 442170 531902 442226
rect 531474 442046 531530 442102
rect 531598 442046 531654 442102
rect 531722 442046 531778 442102
rect 531846 442046 531902 442102
rect 531474 441922 531530 441978
rect 531598 441922 531654 441978
rect 531722 441922 531778 441978
rect 531846 441922 531902 441978
rect 531474 424294 531530 424350
rect 531598 424294 531654 424350
rect 531722 424294 531778 424350
rect 531846 424294 531902 424350
rect 531474 424170 531530 424226
rect 531598 424170 531654 424226
rect 531722 424170 531778 424226
rect 531846 424170 531902 424226
rect 531474 424046 531530 424102
rect 531598 424046 531654 424102
rect 531722 424046 531778 424102
rect 531846 424046 531902 424102
rect 531474 423922 531530 423978
rect 531598 423922 531654 423978
rect 531722 423922 531778 423978
rect 531846 423922 531902 423978
rect 531474 406294 531530 406350
rect 531598 406294 531654 406350
rect 531722 406294 531778 406350
rect 531846 406294 531902 406350
rect 531474 406170 531530 406226
rect 531598 406170 531654 406226
rect 531722 406170 531778 406226
rect 531846 406170 531902 406226
rect 531474 406046 531530 406102
rect 531598 406046 531654 406102
rect 531722 406046 531778 406102
rect 531846 406046 531902 406102
rect 531474 405922 531530 405978
rect 531598 405922 531654 405978
rect 531722 405922 531778 405978
rect 531846 405922 531902 405978
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 551318 514294 551374 514350
rect 551442 514294 551498 514350
rect 551318 514170 551374 514226
rect 551442 514170 551498 514226
rect 551318 514046 551374 514102
rect 551442 514046 551498 514102
rect 551318 513922 551374 513978
rect 551442 513922 551498 513978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 551318 496294 551374 496350
rect 551442 496294 551498 496350
rect 551318 496170 551374 496226
rect 551442 496170 551498 496226
rect 551318 496046 551374 496102
rect 551442 496046 551498 496102
rect 551318 495922 551374 495978
rect 551442 495922 551498 495978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 551318 478294 551374 478350
rect 551442 478294 551498 478350
rect 551318 478170 551374 478226
rect 551442 478170 551498 478226
rect 551318 478046 551374 478102
rect 551442 478046 551498 478102
rect 551318 477922 551374 477978
rect 551442 477922 551498 477978
rect 558474 472294 558530 472350
rect 558598 472294 558654 472350
rect 558722 472294 558778 472350
rect 558846 472294 558902 472350
rect 558474 472170 558530 472226
rect 558598 472170 558654 472226
rect 558722 472170 558778 472226
rect 558846 472170 558902 472226
rect 558474 472046 558530 472102
rect 558598 472046 558654 472102
rect 558722 472046 558778 472102
rect 558846 472046 558902 472102
rect 558474 471922 558530 471978
rect 558598 471922 558654 471978
rect 558722 471922 558778 471978
rect 558846 471922 558902 471978
rect 551318 460294 551374 460350
rect 551442 460294 551498 460350
rect 551318 460170 551374 460226
rect 551442 460170 551498 460226
rect 551318 460046 551374 460102
rect 551442 460046 551498 460102
rect 551318 459922 551374 459978
rect 551442 459922 551498 459978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 558474 400294 558530 400350
rect 558598 400294 558654 400350
rect 558722 400294 558778 400350
rect 558846 400294 558902 400350
rect 558474 400170 558530 400226
rect 558598 400170 558654 400226
rect 558722 400170 558778 400226
rect 558846 400170 558902 400226
rect 558474 400046 558530 400102
rect 558598 400046 558654 400102
rect 558722 400046 558778 400102
rect 558846 400046 558902 400102
rect 558474 399922 558530 399978
rect 558598 399922 558654 399978
rect 558722 399922 558778 399978
rect 558846 399922 558902 399978
rect 531474 388294 531530 388350
rect 531598 388294 531654 388350
rect 531722 388294 531778 388350
rect 531846 388294 531902 388350
rect 531474 388170 531530 388226
rect 531598 388170 531654 388226
rect 531722 388170 531778 388226
rect 531846 388170 531902 388226
rect 531474 388046 531530 388102
rect 531598 388046 531654 388102
rect 531722 388046 531778 388102
rect 531846 388046 531902 388102
rect 531474 387922 531530 387978
rect 531598 387922 531654 387978
rect 531722 387922 531778 387978
rect 531846 387922 531902 387978
rect 531474 370294 531530 370350
rect 531598 370294 531654 370350
rect 531722 370294 531778 370350
rect 531846 370294 531902 370350
rect 531474 370170 531530 370226
rect 531598 370170 531654 370226
rect 531722 370170 531778 370226
rect 531846 370170 531902 370226
rect 531474 370046 531530 370102
rect 531598 370046 531654 370102
rect 531722 370046 531778 370102
rect 531846 370046 531902 370102
rect 531474 369922 531530 369978
rect 531598 369922 531654 369978
rect 531722 369922 531778 369978
rect 531846 369922 531902 369978
rect 531474 352294 531530 352350
rect 531598 352294 531654 352350
rect 531722 352294 531778 352350
rect 531846 352294 531902 352350
rect 531474 352170 531530 352226
rect 531598 352170 531654 352226
rect 531722 352170 531778 352226
rect 531846 352170 531902 352226
rect 531474 352046 531530 352102
rect 531598 352046 531654 352102
rect 531722 352046 531778 352102
rect 531846 352046 531902 352102
rect 531474 351922 531530 351978
rect 531598 351922 531654 351978
rect 531722 351922 531778 351978
rect 531846 351922 531902 351978
rect 531474 334294 531530 334350
rect 531598 334294 531654 334350
rect 531722 334294 531778 334350
rect 531846 334294 531902 334350
rect 531474 334170 531530 334226
rect 531598 334170 531654 334226
rect 531722 334170 531778 334226
rect 531846 334170 531902 334226
rect 531474 334046 531530 334102
rect 531598 334046 531654 334102
rect 531722 334046 531778 334102
rect 531846 334046 531902 334102
rect 531474 333922 531530 333978
rect 531598 333922 531654 333978
rect 531722 333922 531778 333978
rect 531846 333922 531902 333978
rect 531474 316294 531530 316350
rect 531598 316294 531654 316350
rect 531722 316294 531778 316350
rect 531846 316294 531902 316350
rect 531474 316170 531530 316226
rect 531598 316170 531654 316226
rect 531722 316170 531778 316226
rect 531846 316170 531902 316226
rect 531474 316046 531530 316102
rect 531598 316046 531654 316102
rect 531722 316046 531778 316102
rect 531846 316046 531902 316102
rect 531474 315922 531530 315978
rect 531598 315922 531654 315978
rect 531722 315922 531778 315978
rect 531846 315922 531902 315978
rect 531474 298294 531530 298350
rect 531598 298294 531654 298350
rect 531722 298294 531778 298350
rect 531846 298294 531902 298350
rect 531474 298170 531530 298226
rect 531598 298170 531654 298226
rect 531722 298170 531778 298226
rect 531846 298170 531902 298226
rect 531474 298046 531530 298102
rect 531598 298046 531654 298102
rect 531722 298046 531778 298102
rect 531846 298046 531902 298102
rect 531474 297922 531530 297978
rect 531598 297922 531654 297978
rect 531722 297922 531778 297978
rect 531846 297922 531902 297978
rect 531474 280294 531530 280350
rect 531598 280294 531654 280350
rect 531722 280294 531778 280350
rect 531846 280294 531902 280350
rect 531474 280170 531530 280226
rect 531598 280170 531654 280226
rect 531722 280170 531778 280226
rect 531846 280170 531902 280226
rect 531474 280046 531530 280102
rect 531598 280046 531654 280102
rect 531722 280046 531778 280102
rect 531846 280046 531902 280102
rect 531474 279922 531530 279978
rect 531598 279922 531654 279978
rect 531722 279922 531778 279978
rect 531846 279922 531902 279978
rect 531474 262294 531530 262350
rect 531598 262294 531654 262350
rect 531722 262294 531778 262350
rect 531846 262294 531902 262350
rect 531474 262170 531530 262226
rect 531598 262170 531654 262226
rect 531722 262170 531778 262226
rect 531846 262170 531902 262226
rect 531474 262046 531530 262102
rect 531598 262046 531654 262102
rect 531722 262046 531778 262102
rect 531846 262046 531902 262102
rect 531474 261922 531530 261978
rect 531598 261922 531654 261978
rect 531722 261922 531778 261978
rect 531846 261922 531902 261978
rect 558474 382294 558530 382350
rect 558598 382294 558654 382350
rect 558722 382294 558778 382350
rect 558846 382294 558902 382350
rect 558474 382170 558530 382226
rect 558598 382170 558654 382226
rect 558722 382170 558778 382226
rect 558846 382170 558902 382226
rect 558474 382046 558530 382102
rect 558598 382046 558654 382102
rect 558722 382046 558778 382102
rect 558846 382046 558902 382102
rect 558474 381922 558530 381978
rect 558598 381922 558654 381978
rect 558722 381922 558778 381978
rect 558846 381922 558902 381978
rect 558474 364294 558530 364350
rect 558598 364294 558654 364350
rect 558722 364294 558778 364350
rect 558846 364294 558902 364350
rect 558474 364170 558530 364226
rect 558598 364170 558654 364226
rect 558722 364170 558778 364226
rect 558846 364170 558902 364226
rect 558474 364046 558530 364102
rect 558598 364046 558654 364102
rect 558722 364046 558778 364102
rect 558846 364046 558902 364102
rect 558474 363922 558530 363978
rect 558598 363922 558654 363978
rect 558722 363922 558778 363978
rect 558846 363922 558902 363978
rect 558474 346294 558530 346350
rect 558598 346294 558654 346350
rect 558722 346294 558778 346350
rect 558846 346294 558902 346350
rect 558474 346170 558530 346226
rect 558598 346170 558654 346226
rect 558722 346170 558778 346226
rect 558846 346170 558902 346226
rect 558474 346046 558530 346102
rect 558598 346046 558654 346102
rect 558722 346046 558778 346102
rect 558846 346046 558902 346102
rect 558474 345922 558530 345978
rect 558598 345922 558654 345978
rect 558722 345922 558778 345978
rect 558846 345922 558902 345978
rect 558474 328294 558530 328350
rect 558598 328294 558654 328350
rect 558722 328294 558778 328350
rect 558846 328294 558902 328350
rect 558474 328170 558530 328226
rect 558598 328170 558654 328226
rect 558722 328170 558778 328226
rect 558846 328170 558902 328226
rect 558474 328046 558530 328102
rect 558598 328046 558654 328102
rect 558722 328046 558778 328102
rect 558846 328046 558902 328102
rect 558474 327922 558530 327978
rect 558598 327922 558654 327978
rect 558722 327922 558778 327978
rect 558846 327922 558902 327978
rect 558474 310294 558530 310350
rect 558598 310294 558654 310350
rect 558722 310294 558778 310350
rect 558846 310294 558902 310350
rect 558474 310170 558530 310226
rect 558598 310170 558654 310226
rect 558722 310170 558778 310226
rect 558846 310170 558902 310226
rect 558474 310046 558530 310102
rect 558598 310046 558654 310102
rect 558722 310046 558778 310102
rect 558846 310046 558902 310102
rect 558474 309922 558530 309978
rect 558598 309922 558654 309978
rect 558722 309922 558778 309978
rect 558846 309922 558902 309978
rect 558474 292294 558530 292350
rect 558598 292294 558654 292350
rect 558722 292294 558778 292350
rect 558846 292294 558902 292350
rect 558474 292170 558530 292226
rect 558598 292170 558654 292226
rect 558722 292170 558778 292226
rect 558846 292170 558902 292226
rect 558474 292046 558530 292102
rect 558598 292046 558654 292102
rect 558722 292046 558778 292102
rect 558846 292046 558902 292102
rect 558474 291922 558530 291978
rect 558598 291922 558654 291978
rect 558722 291922 558778 291978
rect 558846 291922 558902 291978
rect 558474 274294 558530 274350
rect 558598 274294 558654 274350
rect 558722 274294 558778 274350
rect 558846 274294 558902 274350
rect 558474 274170 558530 274226
rect 558598 274170 558654 274226
rect 558722 274170 558778 274226
rect 558846 274170 558902 274226
rect 558474 274046 558530 274102
rect 558598 274046 558654 274102
rect 558722 274046 558778 274102
rect 558846 274046 558902 274102
rect 558474 273922 558530 273978
rect 558598 273922 558654 273978
rect 558722 273922 558778 273978
rect 558846 273922 558902 273978
rect 558474 256294 558530 256350
rect 558598 256294 558654 256350
rect 558722 256294 558778 256350
rect 558846 256294 558902 256350
rect 558474 256170 558530 256226
rect 558598 256170 558654 256226
rect 558722 256170 558778 256226
rect 558846 256170 558902 256226
rect 558474 256046 558530 256102
rect 558598 256046 558654 256102
rect 558722 256046 558778 256102
rect 558846 256046 558902 256102
rect 557414 255967 557470 256023
rect 557538 255967 557594 256023
rect 557662 255967 557718 256023
rect 557786 255967 557842 256023
rect 557414 255843 557470 255899
rect 557538 255843 557594 255899
rect 557662 255843 557718 255899
rect 557786 255843 557842 255899
rect 558474 255922 558530 255978
rect 558598 255922 558654 255978
rect 558722 255922 558778 255978
rect 558846 255922 558902 255978
rect 531474 244294 531530 244350
rect 531598 244294 531654 244350
rect 531722 244294 531778 244350
rect 531846 244294 531902 244350
rect 531474 244170 531530 244226
rect 531598 244170 531654 244226
rect 531722 244170 531778 244226
rect 531846 244170 531902 244226
rect 531474 244046 531530 244102
rect 531598 244046 531654 244102
rect 531722 244046 531778 244102
rect 531846 244046 531902 244102
rect 531474 243922 531530 243978
rect 531598 243922 531654 243978
rect 531722 243922 531778 243978
rect 531846 243922 531902 243978
rect 556614 244294 556670 244350
rect 556738 244294 556794 244350
rect 556862 244294 556918 244350
rect 556986 244294 557042 244350
rect 556614 244170 556670 244226
rect 556738 244170 556794 244226
rect 556862 244170 556918 244226
rect 556986 244170 557042 244226
rect 556614 244046 556670 244102
rect 556738 244046 556794 244102
rect 556862 244046 556918 244102
rect 556986 244046 557042 244102
rect 556614 243922 556670 243978
rect 556738 243922 556794 243978
rect 556862 243922 556918 243978
rect 556986 243922 557042 243978
rect 557414 238294 557470 238350
rect 557538 238294 557594 238350
rect 557662 238294 557718 238350
rect 557786 238294 557842 238350
rect 557414 238170 557470 238226
rect 557538 238170 557594 238226
rect 557662 238170 557718 238226
rect 557786 238170 557842 238226
rect 557414 238046 557470 238102
rect 557538 238046 557594 238102
rect 557662 238046 557718 238102
rect 557786 238046 557842 238102
rect 557414 237922 557470 237978
rect 557538 237922 557594 237978
rect 557662 237922 557718 237978
rect 557786 237922 557842 237978
rect 558474 238294 558530 238350
rect 558598 238294 558654 238350
rect 558722 238294 558778 238350
rect 558846 238294 558902 238350
rect 558474 238170 558530 238226
rect 558598 238170 558654 238226
rect 558722 238170 558778 238226
rect 558846 238170 558902 238226
rect 558474 238046 558530 238102
rect 558598 238046 558654 238102
rect 558722 238046 558778 238102
rect 558846 238046 558902 238102
rect 558474 237922 558530 237978
rect 558598 237922 558654 237978
rect 558722 237922 558778 237978
rect 558846 237922 558902 237978
rect 531474 226294 531530 226350
rect 531598 226294 531654 226350
rect 531722 226294 531778 226350
rect 531846 226294 531902 226350
rect 531474 226170 531530 226226
rect 531598 226170 531654 226226
rect 531722 226170 531778 226226
rect 531846 226170 531902 226226
rect 531474 226046 531530 226102
rect 531598 226046 531654 226102
rect 531722 226046 531778 226102
rect 531846 226046 531902 226102
rect 531474 225922 531530 225978
rect 531598 225922 531654 225978
rect 531722 225922 531778 225978
rect 531846 225922 531902 225978
rect 556614 226294 556670 226350
rect 556738 226294 556794 226350
rect 556862 226294 556918 226350
rect 556986 226294 557042 226350
rect 556614 226170 556670 226226
rect 556738 226170 556794 226226
rect 556862 226170 556918 226226
rect 556986 226170 557042 226226
rect 556614 226046 556670 226102
rect 556738 226046 556794 226102
rect 556862 226046 556918 226102
rect 556986 226046 557042 226102
rect 556614 225922 556670 225978
rect 556738 225922 556794 225978
rect 556862 225922 556918 225978
rect 556986 225922 557042 225978
rect 557414 220294 557470 220350
rect 557538 220294 557594 220350
rect 557662 220294 557718 220350
rect 557786 220294 557842 220350
rect 557414 220170 557470 220226
rect 557538 220170 557594 220226
rect 557662 220170 557718 220226
rect 557786 220170 557842 220226
rect 557414 220046 557470 220102
rect 557538 220046 557594 220102
rect 557662 220046 557718 220102
rect 557786 220046 557842 220102
rect 557414 219922 557470 219978
rect 557538 219922 557594 219978
rect 557662 219922 557718 219978
rect 557786 219922 557842 219978
rect 558474 220294 558530 220350
rect 558598 220294 558654 220350
rect 558722 220294 558778 220350
rect 558846 220294 558902 220350
rect 558474 220170 558530 220226
rect 558598 220170 558654 220226
rect 558722 220170 558778 220226
rect 558846 220170 558902 220226
rect 558474 220046 558530 220102
rect 558598 220046 558654 220102
rect 558722 220046 558778 220102
rect 558846 220046 558902 220102
rect 558474 219922 558530 219978
rect 558598 219922 558654 219978
rect 558722 219922 558778 219978
rect 558846 219922 558902 219978
rect 531474 208294 531530 208350
rect 531598 208294 531654 208350
rect 531722 208294 531778 208350
rect 531846 208294 531902 208350
rect 531474 208170 531530 208226
rect 531598 208170 531654 208226
rect 531722 208170 531778 208226
rect 531846 208170 531902 208226
rect 531474 208046 531530 208102
rect 531598 208046 531654 208102
rect 531722 208046 531778 208102
rect 531846 208046 531902 208102
rect 531474 207922 531530 207978
rect 531598 207922 531654 207978
rect 531722 207922 531778 207978
rect 531846 207922 531902 207978
rect 556614 208294 556670 208350
rect 556738 208294 556794 208350
rect 556862 208294 556918 208350
rect 556986 208294 557042 208350
rect 556614 208170 556670 208226
rect 556738 208170 556794 208226
rect 556862 208170 556918 208226
rect 556986 208170 557042 208226
rect 556614 208046 556670 208102
rect 556738 208046 556794 208102
rect 556862 208046 556918 208102
rect 556986 208046 557042 208102
rect 556614 207922 556670 207978
rect 556738 207922 556794 207978
rect 556862 207922 556918 207978
rect 556986 207922 557042 207978
rect 557414 202294 557470 202350
rect 557538 202294 557594 202350
rect 557662 202294 557718 202350
rect 557786 202294 557842 202350
rect 557414 202170 557470 202226
rect 557538 202170 557594 202226
rect 557662 202170 557718 202226
rect 557786 202170 557842 202226
rect 557414 202046 557470 202102
rect 557538 202046 557594 202102
rect 557662 202046 557718 202102
rect 557786 202046 557842 202102
rect 557414 201922 557470 201978
rect 557538 201922 557594 201978
rect 557662 201922 557718 201978
rect 557786 201922 557842 201978
rect 558474 202294 558530 202350
rect 558598 202294 558654 202350
rect 558722 202294 558778 202350
rect 558846 202294 558902 202350
rect 558474 202170 558530 202226
rect 558598 202170 558654 202226
rect 558722 202170 558778 202226
rect 558846 202170 558902 202226
rect 558474 202046 558530 202102
rect 558598 202046 558654 202102
rect 558722 202046 558778 202102
rect 558846 202046 558902 202102
rect 558474 201922 558530 201978
rect 558598 201922 558654 201978
rect 558722 201922 558778 201978
rect 558846 201922 558902 201978
rect 531474 190294 531530 190350
rect 531598 190294 531654 190350
rect 531722 190294 531778 190350
rect 531846 190294 531902 190350
rect 531474 190170 531530 190226
rect 531598 190170 531654 190226
rect 531722 190170 531778 190226
rect 531846 190170 531902 190226
rect 531474 190046 531530 190102
rect 531598 190046 531654 190102
rect 531722 190046 531778 190102
rect 531846 190046 531902 190102
rect 531474 189922 531530 189978
rect 531598 189922 531654 189978
rect 531722 189922 531778 189978
rect 531846 189922 531902 189978
rect 556614 190294 556670 190350
rect 556738 190294 556794 190350
rect 556862 190294 556918 190350
rect 556986 190294 557042 190350
rect 556614 190170 556670 190226
rect 556738 190170 556794 190226
rect 556862 190170 556918 190226
rect 556986 190170 557042 190226
rect 556614 190046 556670 190102
rect 556738 190046 556794 190102
rect 556862 190046 556918 190102
rect 556986 190046 557042 190102
rect 556614 189922 556670 189978
rect 556738 189922 556794 189978
rect 556862 189922 556918 189978
rect 556986 189922 557042 189978
rect 557414 184294 557470 184350
rect 557538 184294 557594 184350
rect 557662 184294 557718 184350
rect 557786 184294 557842 184350
rect 557414 184170 557470 184226
rect 557538 184170 557594 184226
rect 557662 184170 557718 184226
rect 557786 184170 557842 184226
rect 557414 184046 557470 184102
rect 557538 184046 557594 184102
rect 557662 184046 557718 184102
rect 557786 184046 557842 184102
rect 557414 183922 557470 183978
rect 557538 183922 557594 183978
rect 557662 183922 557718 183978
rect 557786 183922 557842 183978
rect 558474 184294 558530 184350
rect 558598 184294 558654 184350
rect 558722 184294 558778 184350
rect 558846 184294 558902 184350
rect 558474 184170 558530 184226
rect 558598 184170 558654 184226
rect 558722 184170 558778 184226
rect 558846 184170 558902 184226
rect 558474 184046 558530 184102
rect 558598 184046 558654 184102
rect 558722 184046 558778 184102
rect 558846 184046 558902 184102
rect 558474 183922 558530 183978
rect 558598 183922 558654 183978
rect 558722 183922 558778 183978
rect 558846 183922 558902 183978
rect 531474 172294 531530 172350
rect 531598 172294 531654 172350
rect 531722 172294 531778 172350
rect 531846 172294 531902 172350
rect 531474 172170 531530 172226
rect 531598 172170 531654 172226
rect 531722 172170 531778 172226
rect 531846 172170 531902 172226
rect 531474 172046 531530 172102
rect 531598 172046 531654 172102
rect 531722 172046 531778 172102
rect 531846 172046 531902 172102
rect 531474 171922 531530 171978
rect 531598 171922 531654 171978
rect 531722 171922 531778 171978
rect 531846 171922 531902 171978
rect 556614 172294 556670 172350
rect 556738 172294 556794 172350
rect 556862 172294 556918 172350
rect 556986 172294 557042 172350
rect 556614 172170 556670 172226
rect 556738 172170 556794 172226
rect 556862 172170 556918 172226
rect 556986 172170 557042 172226
rect 556614 172046 556670 172102
rect 556738 172046 556794 172102
rect 556862 172046 556918 172102
rect 556986 172046 557042 172102
rect 556614 171922 556670 171978
rect 556738 171922 556794 171978
rect 556862 171922 556918 171978
rect 556986 171922 557042 171978
rect 557414 166294 557470 166350
rect 557538 166294 557594 166350
rect 557662 166294 557718 166350
rect 557786 166294 557842 166350
rect 557414 166170 557470 166226
rect 557538 166170 557594 166226
rect 557662 166170 557718 166226
rect 557786 166170 557842 166226
rect 557414 166046 557470 166102
rect 557538 166046 557594 166102
rect 557662 166046 557718 166102
rect 557786 166046 557842 166102
rect 557414 165922 557470 165978
rect 557538 165922 557594 165978
rect 557662 165922 557718 165978
rect 557786 165922 557842 165978
rect 558474 166294 558530 166350
rect 558598 166294 558654 166350
rect 558722 166294 558778 166350
rect 558846 166294 558902 166350
rect 558474 166170 558530 166226
rect 558598 166170 558654 166226
rect 558722 166170 558778 166226
rect 558846 166170 558902 166226
rect 558474 166046 558530 166102
rect 558598 166046 558654 166102
rect 558722 166046 558778 166102
rect 558846 166046 558902 166102
rect 558474 165922 558530 165978
rect 558598 165922 558654 165978
rect 558722 165922 558778 165978
rect 558846 165922 558902 165978
rect 531474 154294 531530 154350
rect 531598 154294 531654 154350
rect 531722 154294 531778 154350
rect 531846 154294 531902 154350
rect 531474 154170 531530 154226
rect 531598 154170 531654 154226
rect 531722 154170 531778 154226
rect 531846 154170 531902 154226
rect 531474 154046 531530 154102
rect 531598 154046 531654 154102
rect 531722 154046 531778 154102
rect 531846 154046 531902 154102
rect 531474 153922 531530 153978
rect 531598 153922 531654 153978
rect 531722 153922 531778 153978
rect 531846 153922 531902 153978
rect 558474 148294 558530 148350
rect 558598 148294 558654 148350
rect 558722 148294 558778 148350
rect 558846 148294 558902 148350
rect 558474 148170 558530 148226
rect 558598 148170 558654 148226
rect 558722 148170 558778 148226
rect 558846 148170 558902 148226
rect 558474 148046 558530 148102
rect 558598 148046 558654 148102
rect 558722 148046 558778 148102
rect 558846 148046 558902 148102
rect 558474 147922 558530 147978
rect 558598 147922 558654 147978
rect 558722 147922 558778 147978
rect 558846 147922 558902 147978
rect 544684 142442 544740 142498
rect 534604 141902 534660 141958
rect 531474 136294 531530 136350
rect 531598 136294 531654 136350
rect 531722 136294 531778 136350
rect 531846 136294 531902 136350
rect 531474 136170 531530 136226
rect 531598 136170 531654 136226
rect 531722 136170 531778 136226
rect 531846 136170 531902 136226
rect 531474 136046 531530 136102
rect 531598 136046 531654 136102
rect 531722 136046 531778 136102
rect 531846 136046 531902 136102
rect 531474 135922 531530 135978
rect 531598 135922 531654 135978
rect 531722 135922 531778 135978
rect 531846 135922 531902 135978
rect 545812 130294 545868 130350
rect 545936 130294 545992 130350
rect 546060 130294 546116 130350
rect 546184 130294 546240 130350
rect 545812 130170 545868 130226
rect 545936 130170 545992 130226
rect 546060 130170 546116 130226
rect 546184 130170 546240 130226
rect 545812 130046 545868 130102
rect 545936 130046 545992 130102
rect 546060 130046 546116 130102
rect 546184 130046 546240 130102
rect 545812 129922 545868 129978
rect 545936 129922 545992 129978
rect 546060 129922 546116 129978
rect 546184 129922 546240 129978
rect 558474 130294 558530 130350
rect 558598 130294 558654 130350
rect 558722 130294 558778 130350
rect 558846 130294 558902 130350
rect 558474 130170 558530 130226
rect 558598 130170 558654 130226
rect 558722 130170 558778 130226
rect 558846 130170 558902 130226
rect 558474 130046 558530 130102
rect 558598 130046 558654 130102
rect 558722 130046 558778 130102
rect 558846 130046 558902 130102
rect 558474 129922 558530 129978
rect 558598 129922 558654 129978
rect 558722 129922 558778 129978
rect 558846 129922 558902 129978
rect 531474 118294 531530 118350
rect 531598 118294 531654 118350
rect 531722 118294 531778 118350
rect 531846 118294 531902 118350
rect 531474 118170 531530 118226
rect 531598 118170 531654 118226
rect 531722 118170 531778 118226
rect 531846 118170 531902 118226
rect 531474 118046 531530 118102
rect 531598 118046 531654 118102
rect 531722 118046 531778 118102
rect 531846 118046 531902 118102
rect 531474 117922 531530 117978
rect 531598 117922 531654 117978
rect 531722 117922 531778 117978
rect 531846 117922 531902 117978
rect 546612 118294 546668 118350
rect 546736 118294 546792 118350
rect 546860 118294 546916 118350
rect 546984 118294 547040 118350
rect 546612 118170 546668 118226
rect 546736 118170 546792 118226
rect 546860 118170 546916 118226
rect 546984 118170 547040 118226
rect 546612 118046 546668 118102
rect 546736 118046 546792 118102
rect 546860 118046 546916 118102
rect 546984 118046 547040 118102
rect 546612 117922 546668 117978
rect 546736 117922 546792 117978
rect 546860 117922 546916 117978
rect 546984 117922 547040 117978
rect 545812 112294 545868 112350
rect 545936 112294 545992 112350
rect 546060 112294 546116 112350
rect 546184 112294 546240 112350
rect 545812 112170 545868 112226
rect 545936 112170 545992 112226
rect 546060 112170 546116 112226
rect 546184 112170 546240 112226
rect 545812 112046 545868 112102
rect 545936 112046 545992 112102
rect 546060 112046 546116 112102
rect 546184 112046 546240 112102
rect 545812 111922 545868 111978
rect 545936 111922 545992 111978
rect 546060 111922 546116 111978
rect 546184 111922 546240 111978
rect 558474 112294 558530 112350
rect 558598 112294 558654 112350
rect 558722 112294 558778 112350
rect 558846 112294 558902 112350
rect 558474 112170 558530 112226
rect 558598 112170 558654 112226
rect 558722 112170 558778 112226
rect 558846 112170 558902 112226
rect 558474 112046 558530 112102
rect 558598 112046 558654 112102
rect 558722 112046 558778 112102
rect 558846 112046 558902 112102
rect 558474 111922 558530 111978
rect 558598 111922 558654 111978
rect 558722 111922 558778 111978
rect 558846 111922 558902 111978
rect 531474 100294 531530 100350
rect 531598 100294 531654 100350
rect 531722 100294 531778 100350
rect 531846 100294 531902 100350
rect 531474 100170 531530 100226
rect 531598 100170 531654 100226
rect 531722 100170 531778 100226
rect 531846 100170 531902 100226
rect 531474 100046 531530 100102
rect 531598 100046 531654 100102
rect 531722 100046 531778 100102
rect 531846 100046 531902 100102
rect 531474 99922 531530 99978
rect 531598 99922 531654 99978
rect 531722 99922 531778 99978
rect 531846 99922 531902 99978
rect 546612 100294 546668 100350
rect 546736 100294 546792 100350
rect 546860 100294 546916 100350
rect 546984 100294 547040 100350
rect 546612 100170 546668 100226
rect 546736 100170 546792 100226
rect 546860 100170 546916 100226
rect 546984 100170 547040 100226
rect 546612 100046 546668 100102
rect 546736 100046 546792 100102
rect 546860 100046 546916 100102
rect 546984 100046 547040 100102
rect 546612 99922 546668 99978
rect 546736 99922 546792 99978
rect 546860 99922 546916 99978
rect 546984 99922 547040 99978
rect 545812 94294 545868 94350
rect 545936 94294 545992 94350
rect 546060 94294 546116 94350
rect 546184 94294 546240 94350
rect 545812 94170 545868 94226
rect 545936 94170 545992 94226
rect 546060 94170 546116 94226
rect 546184 94170 546240 94226
rect 545812 94046 545868 94102
rect 545936 94046 545992 94102
rect 546060 94046 546116 94102
rect 546184 94046 546240 94102
rect 545812 93922 545868 93978
rect 545936 93922 545992 93978
rect 546060 93922 546116 93978
rect 546184 93922 546240 93978
rect 558474 94294 558530 94350
rect 558598 94294 558654 94350
rect 558722 94294 558778 94350
rect 558846 94294 558902 94350
rect 558474 94170 558530 94226
rect 558598 94170 558654 94226
rect 558722 94170 558778 94226
rect 558846 94170 558902 94226
rect 558474 94046 558530 94102
rect 558598 94046 558654 94102
rect 558722 94046 558778 94102
rect 558846 94046 558902 94102
rect 558474 93922 558530 93978
rect 558598 93922 558654 93978
rect 558722 93922 558778 93978
rect 558846 93922 558902 93978
rect 531474 82294 531530 82350
rect 531598 82294 531654 82350
rect 531722 82294 531778 82350
rect 531846 82294 531902 82350
rect 531474 82170 531530 82226
rect 531598 82170 531654 82226
rect 531722 82170 531778 82226
rect 531846 82170 531902 82226
rect 531474 82046 531530 82102
rect 531598 82046 531654 82102
rect 531722 82046 531778 82102
rect 531846 82046 531902 82102
rect 531474 81922 531530 81978
rect 531598 81922 531654 81978
rect 531722 81922 531778 81978
rect 531846 81922 531902 81978
rect 546612 82294 546668 82350
rect 546736 82294 546792 82350
rect 546860 82294 546916 82350
rect 546984 82294 547040 82350
rect 546612 82170 546668 82226
rect 546736 82170 546792 82226
rect 546860 82170 546916 82226
rect 546984 82170 547040 82226
rect 546612 82046 546668 82102
rect 546736 82046 546792 82102
rect 546860 82046 546916 82102
rect 546984 82046 547040 82102
rect 546612 81922 546668 81978
rect 546736 81922 546792 81978
rect 546860 81922 546916 81978
rect 546984 81922 547040 81978
rect 545812 76294 545868 76350
rect 545936 76294 545992 76350
rect 546060 76294 546116 76350
rect 546184 76294 546240 76350
rect 545812 76170 545868 76226
rect 545936 76170 545992 76226
rect 546060 76170 546116 76226
rect 546184 76170 546240 76226
rect 545812 76046 545868 76102
rect 545936 76046 545992 76102
rect 546060 76046 546116 76102
rect 546184 76046 546240 76102
rect 545812 75922 545868 75978
rect 545936 75922 545992 75978
rect 546060 75922 546116 75978
rect 546184 75922 546240 75978
rect 558474 76294 558530 76350
rect 558598 76294 558654 76350
rect 558722 76294 558778 76350
rect 558846 76294 558902 76350
rect 558474 76170 558530 76226
rect 558598 76170 558654 76226
rect 558722 76170 558778 76226
rect 558846 76170 558902 76226
rect 558474 76046 558530 76102
rect 558598 76046 558654 76102
rect 558722 76046 558778 76102
rect 558846 76046 558902 76102
rect 558474 75922 558530 75978
rect 558598 75922 558654 75978
rect 558722 75922 558778 75978
rect 558846 75922 558902 75978
rect 531474 64294 531530 64350
rect 531598 64294 531654 64350
rect 531722 64294 531778 64350
rect 531846 64294 531902 64350
rect 531474 64170 531530 64226
rect 531598 64170 531654 64226
rect 531722 64170 531778 64226
rect 531846 64170 531902 64226
rect 531474 64046 531530 64102
rect 531598 64046 531654 64102
rect 531722 64046 531778 64102
rect 531846 64046 531902 64102
rect 531474 63922 531530 63978
rect 531598 63922 531654 63978
rect 531722 63922 531778 63978
rect 531846 63922 531902 63978
rect 546612 64294 546668 64350
rect 546736 64294 546792 64350
rect 546860 64294 546916 64350
rect 546984 64294 547040 64350
rect 546612 64170 546668 64226
rect 546736 64170 546792 64226
rect 546860 64170 546916 64226
rect 546984 64170 547040 64226
rect 546612 64046 546668 64102
rect 546736 64046 546792 64102
rect 546860 64046 546916 64102
rect 546984 64046 547040 64102
rect 546612 63922 546668 63978
rect 546736 63922 546792 63978
rect 546860 63922 546916 63978
rect 546984 63922 547040 63978
rect 545812 58294 545868 58350
rect 545936 58294 545992 58350
rect 546060 58294 546116 58350
rect 546184 58294 546240 58350
rect 545812 58170 545868 58226
rect 545936 58170 545992 58226
rect 546060 58170 546116 58226
rect 546184 58170 546240 58226
rect 545812 58046 545868 58102
rect 545936 58046 545992 58102
rect 546060 58046 546116 58102
rect 546184 58046 546240 58102
rect 545812 57922 545868 57978
rect 545936 57922 545992 57978
rect 546060 57922 546116 57978
rect 546184 57922 546240 57978
rect 558474 58294 558530 58350
rect 558598 58294 558654 58350
rect 558722 58294 558778 58350
rect 558846 58294 558902 58350
rect 558474 58170 558530 58226
rect 558598 58170 558654 58226
rect 558722 58170 558778 58226
rect 558846 58170 558902 58226
rect 558474 58046 558530 58102
rect 558598 58046 558654 58102
rect 558722 58046 558778 58102
rect 558846 58046 558902 58102
rect 558474 57922 558530 57978
rect 558598 57922 558654 57978
rect 558722 57922 558778 57978
rect 558846 57922 558902 57978
rect 531474 46294 531530 46350
rect 531598 46294 531654 46350
rect 531722 46294 531778 46350
rect 531846 46294 531902 46350
rect 531474 46170 531530 46226
rect 531598 46170 531654 46226
rect 531722 46170 531778 46226
rect 531846 46170 531902 46226
rect 531474 46046 531530 46102
rect 531598 46046 531654 46102
rect 531722 46046 531778 46102
rect 531846 46046 531902 46102
rect 531474 45922 531530 45978
rect 531598 45922 531654 45978
rect 531722 45922 531778 45978
rect 531846 45922 531902 45978
rect 546612 46294 546668 46350
rect 546736 46294 546792 46350
rect 546860 46294 546916 46350
rect 546984 46294 547040 46350
rect 546612 46170 546668 46226
rect 546736 46170 546792 46226
rect 546860 46170 546916 46226
rect 546984 46170 547040 46226
rect 546612 46046 546668 46102
rect 546736 46046 546792 46102
rect 546860 46046 546916 46102
rect 546984 46046 547040 46102
rect 546612 45922 546668 45978
rect 546736 45922 546792 45978
rect 546860 45922 546916 45978
rect 546984 45922 547040 45978
rect 531474 28294 531530 28350
rect 531598 28294 531654 28350
rect 531722 28294 531778 28350
rect 531846 28294 531902 28350
rect 531474 28170 531530 28226
rect 531598 28170 531654 28226
rect 531722 28170 531778 28226
rect 531846 28170 531902 28226
rect 531474 28046 531530 28102
rect 531598 28046 531654 28102
rect 531722 28046 531778 28102
rect 531846 28046 531902 28102
rect 531474 27922 531530 27978
rect 531598 27922 531654 27978
rect 531722 27922 531778 27978
rect 531846 27922 531902 27978
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 558474 40294 558530 40350
rect 558598 40294 558654 40350
rect 558722 40294 558778 40350
rect 558846 40294 558902 40350
rect 558474 40170 558530 40226
rect 558598 40170 558654 40226
rect 558722 40170 558778 40226
rect 558846 40170 558902 40226
rect 558474 40046 558530 40102
rect 558598 40046 558654 40102
rect 558722 40046 558778 40102
rect 558846 40046 558902 40102
rect 558474 39922 558530 39978
rect 558598 39922 558654 39978
rect 558722 39922 558778 39978
rect 558846 39922 558902 39978
rect 558474 22294 558530 22350
rect 558598 22294 558654 22350
rect 558722 22294 558778 22350
rect 558846 22294 558902 22350
rect 558474 22170 558530 22226
rect 558598 22170 558654 22226
rect 558722 22170 558778 22226
rect 558846 22170 558902 22226
rect 558474 22046 558530 22102
rect 558598 22046 558654 22102
rect 558722 22046 558778 22102
rect 558846 22046 558902 22102
rect 558474 21922 558530 21978
rect 558598 21922 558654 21978
rect 558722 21922 558778 21978
rect 558846 21922 558902 21978
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 584668 589742 584724 589798
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 562194 388294 562250 388350
rect 562318 388294 562374 388350
rect 562442 388294 562498 388350
rect 562566 388294 562622 388350
rect 562194 388170 562250 388226
rect 562318 388170 562374 388226
rect 562442 388170 562498 388226
rect 562566 388170 562622 388226
rect 562194 388046 562250 388102
rect 562318 388046 562374 388102
rect 562442 388046 562498 388102
rect 562566 388046 562622 388102
rect 562194 387922 562250 387978
rect 562318 387922 562374 387978
rect 562442 387922 562498 387978
rect 562566 387922 562622 387978
rect 562194 370294 562250 370350
rect 562318 370294 562374 370350
rect 562442 370294 562498 370350
rect 562566 370294 562622 370350
rect 562194 370170 562250 370226
rect 562318 370170 562374 370226
rect 562442 370170 562498 370226
rect 562566 370170 562622 370226
rect 562194 370046 562250 370102
rect 562318 370046 562374 370102
rect 562442 370046 562498 370102
rect 562566 370046 562622 370102
rect 562194 369922 562250 369978
rect 562318 369922 562374 369978
rect 562442 369922 562498 369978
rect 562566 369922 562622 369978
rect 562194 352294 562250 352350
rect 562318 352294 562374 352350
rect 562442 352294 562498 352350
rect 562566 352294 562622 352350
rect 562194 352170 562250 352226
rect 562318 352170 562374 352226
rect 562442 352170 562498 352226
rect 562566 352170 562622 352226
rect 562194 352046 562250 352102
rect 562318 352046 562374 352102
rect 562442 352046 562498 352102
rect 562566 352046 562622 352102
rect 562194 351922 562250 351978
rect 562318 351922 562374 351978
rect 562442 351922 562498 351978
rect 562566 351922 562622 351978
rect 562194 334294 562250 334350
rect 562318 334294 562374 334350
rect 562442 334294 562498 334350
rect 562566 334294 562622 334350
rect 562194 334170 562250 334226
rect 562318 334170 562374 334226
rect 562442 334170 562498 334226
rect 562566 334170 562622 334226
rect 562194 334046 562250 334102
rect 562318 334046 562374 334102
rect 562442 334046 562498 334102
rect 562566 334046 562622 334102
rect 562194 333922 562250 333978
rect 562318 333922 562374 333978
rect 562442 333922 562498 333978
rect 562566 333922 562622 333978
rect 562194 316294 562250 316350
rect 562318 316294 562374 316350
rect 562442 316294 562498 316350
rect 562566 316294 562622 316350
rect 562194 316170 562250 316226
rect 562318 316170 562374 316226
rect 562442 316170 562498 316226
rect 562566 316170 562622 316226
rect 562194 316046 562250 316102
rect 562318 316046 562374 316102
rect 562442 316046 562498 316102
rect 562566 316046 562622 316102
rect 562194 315922 562250 315978
rect 562318 315922 562374 315978
rect 562442 315922 562498 315978
rect 562566 315922 562622 315978
rect 562194 298294 562250 298350
rect 562318 298294 562374 298350
rect 562442 298294 562498 298350
rect 562566 298294 562622 298350
rect 562194 298170 562250 298226
rect 562318 298170 562374 298226
rect 562442 298170 562498 298226
rect 562566 298170 562622 298226
rect 562194 298046 562250 298102
rect 562318 298046 562374 298102
rect 562442 298046 562498 298102
rect 562566 298046 562622 298102
rect 562194 297922 562250 297978
rect 562318 297922 562374 297978
rect 562442 297922 562498 297978
rect 562566 297922 562622 297978
rect 562194 280294 562250 280350
rect 562318 280294 562374 280350
rect 562442 280294 562498 280350
rect 562566 280294 562622 280350
rect 562194 280170 562250 280226
rect 562318 280170 562374 280226
rect 562442 280170 562498 280226
rect 562566 280170 562622 280226
rect 562194 280046 562250 280102
rect 562318 280046 562374 280102
rect 562442 280046 562498 280102
rect 562566 280046 562622 280102
rect 562194 279922 562250 279978
rect 562318 279922 562374 279978
rect 562442 279922 562498 279978
rect 562566 279922 562622 279978
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 590604 551042 590660 551098
rect 590156 547802 590212 547858
rect 590492 547982 590548 548038
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 590156 376442 590212 376498
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 590492 295442 590548 295498
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 590156 285182 590212 285238
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 590716 450962 590772 451018
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 590828 301562 590884 301618
rect 591052 387602 591108 387658
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 590940 300662 590996 300718
rect 590716 285542 590772 285598
rect 591052 297242 591108 297298
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 591276 295622 591332 295678
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 591164 288782 591220 288838
rect 590828 282122 590884 282178
rect 590604 281942 590660 281998
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 562194 262294 562250 262350
rect 562318 262294 562374 262350
rect 562442 262294 562498 262350
rect 562566 262294 562622 262350
rect 562194 262170 562250 262226
rect 562318 262170 562374 262226
rect 562442 262170 562498 262226
rect 562566 262170 562622 262226
rect 562194 262046 562250 262102
rect 562318 262046 562374 262102
rect 562442 262046 562498 262102
rect 562566 262046 562622 262102
rect 562194 261922 562250 261978
rect 562318 261922 562374 261978
rect 562442 261922 562498 261978
rect 562566 261922 562622 261978
rect 562194 244294 562250 244350
rect 562318 244294 562374 244350
rect 562442 244294 562498 244350
rect 562566 244294 562622 244350
rect 562194 244170 562250 244226
rect 562318 244170 562374 244226
rect 562442 244170 562498 244226
rect 562566 244170 562622 244226
rect 562194 244046 562250 244102
rect 562318 244046 562374 244102
rect 562442 244046 562498 244102
rect 562566 244046 562622 244102
rect 562194 243922 562250 243978
rect 562318 243922 562374 243978
rect 562442 243922 562498 243978
rect 562566 243922 562622 243978
rect 562194 226294 562250 226350
rect 562318 226294 562374 226350
rect 562442 226294 562498 226350
rect 562566 226294 562622 226350
rect 562194 226170 562250 226226
rect 562318 226170 562374 226226
rect 562442 226170 562498 226226
rect 562566 226170 562622 226226
rect 562194 226046 562250 226102
rect 562318 226046 562374 226102
rect 562442 226046 562498 226102
rect 562566 226046 562622 226102
rect 562194 225922 562250 225978
rect 562318 225922 562374 225978
rect 562442 225922 562498 225978
rect 562566 225922 562622 225978
rect 562194 208294 562250 208350
rect 562318 208294 562374 208350
rect 562442 208294 562498 208350
rect 562566 208294 562622 208350
rect 562194 208170 562250 208226
rect 562318 208170 562374 208226
rect 562442 208170 562498 208226
rect 562566 208170 562622 208226
rect 562194 208046 562250 208102
rect 562318 208046 562374 208102
rect 562442 208046 562498 208102
rect 562566 208046 562622 208102
rect 562194 207922 562250 207978
rect 562318 207922 562374 207978
rect 562442 207922 562498 207978
rect 562566 207922 562622 207978
rect 562194 190294 562250 190350
rect 562318 190294 562374 190350
rect 562442 190294 562498 190350
rect 562566 190294 562622 190350
rect 562194 190170 562250 190226
rect 562318 190170 562374 190226
rect 562442 190170 562498 190226
rect 562566 190170 562622 190226
rect 562194 190046 562250 190102
rect 562318 190046 562374 190102
rect 562442 190046 562498 190102
rect 562566 190046 562622 190102
rect 562194 189922 562250 189978
rect 562318 189922 562374 189978
rect 562442 189922 562498 189978
rect 562566 189922 562622 189978
rect 562194 172294 562250 172350
rect 562318 172294 562374 172350
rect 562442 172294 562498 172350
rect 562566 172294 562622 172350
rect 562194 172170 562250 172226
rect 562318 172170 562374 172226
rect 562442 172170 562498 172226
rect 562566 172170 562622 172226
rect 562194 172046 562250 172102
rect 562318 172046 562374 172102
rect 562442 172046 562498 172102
rect 562566 172046 562622 172102
rect 562194 171922 562250 171978
rect 562318 171922 562374 171978
rect 562442 171922 562498 171978
rect 562566 171922 562622 171978
rect 562194 154294 562250 154350
rect 562318 154294 562374 154350
rect 562442 154294 562498 154350
rect 562566 154294 562622 154350
rect 562194 154170 562250 154226
rect 562318 154170 562374 154226
rect 562442 154170 562498 154226
rect 562566 154170 562622 154226
rect 562194 154046 562250 154102
rect 562318 154046 562374 154102
rect 562442 154046 562498 154102
rect 562566 154046 562622 154102
rect 562194 153922 562250 153978
rect 562318 153922 562374 153978
rect 562442 153922 562498 153978
rect 562566 153922 562622 153978
rect 562194 136294 562250 136350
rect 562318 136294 562374 136350
rect 562442 136294 562498 136350
rect 562566 136294 562622 136350
rect 562194 136170 562250 136226
rect 562318 136170 562374 136226
rect 562442 136170 562498 136226
rect 562566 136170 562622 136226
rect 562194 136046 562250 136102
rect 562318 136046 562374 136102
rect 562442 136046 562498 136102
rect 562566 136046 562622 136102
rect 562194 135922 562250 135978
rect 562318 135922 562374 135978
rect 562442 135922 562498 135978
rect 562566 135922 562622 135978
rect 562194 118294 562250 118350
rect 562318 118294 562374 118350
rect 562442 118294 562498 118350
rect 562566 118294 562622 118350
rect 562194 118170 562250 118226
rect 562318 118170 562374 118226
rect 562442 118170 562498 118226
rect 562566 118170 562622 118226
rect 562194 118046 562250 118102
rect 562318 118046 562374 118102
rect 562442 118046 562498 118102
rect 562566 118046 562622 118102
rect 562194 117922 562250 117978
rect 562318 117922 562374 117978
rect 562442 117922 562498 117978
rect 562566 117922 562622 117978
rect 562194 100294 562250 100350
rect 562318 100294 562374 100350
rect 562442 100294 562498 100350
rect 562566 100294 562622 100350
rect 562194 100170 562250 100226
rect 562318 100170 562374 100226
rect 562442 100170 562498 100226
rect 562566 100170 562622 100226
rect 562194 100046 562250 100102
rect 562318 100046 562374 100102
rect 562442 100046 562498 100102
rect 562566 100046 562622 100102
rect 562194 99922 562250 99978
rect 562318 99922 562374 99978
rect 562442 99922 562498 99978
rect 562566 99922 562622 99978
rect 562194 82294 562250 82350
rect 562318 82294 562374 82350
rect 562442 82294 562498 82350
rect 562566 82294 562622 82350
rect 562194 82170 562250 82226
rect 562318 82170 562374 82226
rect 562442 82170 562498 82226
rect 562566 82170 562622 82226
rect 562194 82046 562250 82102
rect 562318 82046 562374 82102
rect 562442 82046 562498 82102
rect 562566 82046 562622 82102
rect 562194 81922 562250 81978
rect 562318 81922 562374 81978
rect 562442 81922 562498 81978
rect 562566 81922 562622 81978
rect 562194 64294 562250 64350
rect 562318 64294 562374 64350
rect 562442 64294 562498 64350
rect 562566 64294 562622 64350
rect 562194 64170 562250 64226
rect 562318 64170 562374 64226
rect 562442 64170 562498 64226
rect 562566 64170 562622 64226
rect 562194 64046 562250 64102
rect 562318 64046 562374 64102
rect 562442 64046 562498 64102
rect 562566 64046 562622 64102
rect 562194 63922 562250 63978
rect 562318 63922 562374 63978
rect 562442 63922 562498 63978
rect 562566 63922 562622 63978
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 590156 206342 590212 206398
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 590156 127502 590212 127558
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 562194 46294 562250 46350
rect 562318 46294 562374 46350
rect 562442 46294 562498 46350
rect 562566 46294 562622 46350
rect 562194 46170 562250 46226
rect 562318 46170 562374 46226
rect 562442 46170 562498 46226
rect 562566 46170 562622 46226
rect 562194 46046 562250 46102
rect 562318 46046 562374 46102
rect 562442 46046 562498 46102
rect 562566 46046 562622 46102
rect 562194 45922 562250 45978
rect 562318 45922 562374 45978
rect 562442 45922 562498 45978
rect 562566 45922 562622 45978
rect 562194 28294 562250 28350
rect 562318 28294 562374 28350
rect 562442 28294 562498 28350
rect 562566 28294 562622 28350
rect 562194 28170 562250 28226
rect 562318 28170 562374 28226
rect 562442 28170 562498 28226
rect 562566 28170 562622 28226
rect 562194 28046 562250 28102
rect 562318 28046 562374 28102
rect 562442 28046 562498 28102
rect 562566 28046 562622 28102
rect 562194 27922 562250 27978
rect 562318 27922 562374 27978
rect 562442 27922 562498 27978
rect 562566 27922 562622 27978
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect 288076 589798 584740 589814
rect 288076 589742 288092 589798
rect 288148 589742 584668 589798
rect 584724 589742 584740 589798
rect 288076 589726 584740 589742
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 220554 562350
rect 220610 562294 220678 562350
rect 220734 562294 220802 562350
rect 220858 562294 220926 562350
rect 220982 562294 251274 562350
rect 251330 562294 251398 562350
rect 251454 562294 251522 562350
rect 251578 562294 251646 562350
rect 251702 562294 281994 562350
rect 282050 562294 282118 562350
rect 282174 562294 282242 562350
rect 282298 562294 282366 562350
rect 282422 562294 312714 562350
rect 312770 562294 312838 562350
rect 312894 562294 312962 562350
rect 313018 562294 313086 562350
rect 313142 562294 343434 562350
rect 343490 562294 343558 562350
rect 343614 562294 343682 562350
rect 343738 562294 343806 562350
rect 343862 562294 374154 562350
rect 374210 562294 374278 562350
rect 374334 562294 374402 562350
rect 374458 562294 374526 562350
rect 374582 562294 404874 562350
rect 404930 562294 404998 562350
rect 405054 562294 405122 562350
rect 405178 562294 405246 562350
rect 405302 562294 435594 562350
rect 435650 562294 435718 562350
rect 435774 562294 435842 562350
rect 435898 562294 435966 562350
rect 436022 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 220554 562226
rect 220610 562170 220678 562226
rect 220734 562170 220802 562226
rect 220858 562170 220926 562226
rect 220982 562170 251274 562226
rect 251330 562170 251398 562226
rect 251454 562170 251522 562226
rect 251578 562170 251646 562226
rect 251702 562170 281994 562226
rect 282050 562170 282118 562226
rect 282174 562170 282242 562226
rect 282298 562170 282366 562226
rect 282422 562170 312714 562226
rect 312770 562170 312838 562226
rect 312894 562170 312962 562226
rect 313018 562170 313086 562226
rect 313142 562170 343434 562226
rect 343490 562170 343558 562226
rect 343614 562170 343682 562226
rect 343738 562170 343806 562226
rect 343862 562170 374154 562226
rect 374210 562170 374278 562226
rect 374334 562170 374402 562226
rect 374458 562170 374526 562226
rect 374582 562170 404874 562226
rect 404930 562170 404998 562226
rect 405054 562170 405122 562226
rect 405178 562170 405246 562226
rect 405302 562170 435594 562226
rect 435650 562170 435718 562226
rect 435774 562170 435842 562226
rect 435898 562170 435966 562226
rect 436022 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 220554 562102
rect 220610 562046 220678 562102
rect 220734 562046 220802 562102
rect 220858 562046 220926 562102
rect 220982 562046 251274 562102
rect 251330 562046 251398 562102
rect 251454 562046 251522 562102
rect 251578 562046 251646 562102
rect 251702 562046 281994 562102
rect 282050 562046 282118 562102
rect 282174 562046 282242 562102
rect 282298 562046 282366 562102
rect 282422 562046 312714 562102
rect 312770 562046 312838 562102
rect 312894 562046 312962 562102
rect 313018 562046 313086 562102
rect 313142 562046 343434 562102
rect 343490 562046 343558 562102
rect 343614 562046 343682 562102
rect 343738 562046 343806 562102
rect 343862 562046 374154 562102
rect 374210 562046 374278 562102
rect 374334 562046 374402 562102
rect 374458 562046 374526 562102
rect 374582 562046 404874 562102
rect 404930 562046 404998 562102
rect 405054 562046 405122 562102
rect 405178 562046 405246 562102
rect 405302 562046 435594 562102
rect 435650 562046 435718 562102
rect 435774 562046 435842 562102
rect 435898 562046 435966 562102
rect 436022 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 220554 561978
rect 220610 561922 220678 561978
rect 220734 561922 220802 561978
rect 220858 561922 220926 561978
rect 220982 561922 251274 561978
rect 251330 561922 251398 561978
rect 251454 561922 251522 561978
rect 251578 561922 251646 561978
rect 251702 561922 281994 561978
rect 282050 561922 282118 561978
rect 282174 561922 282242 561978
rect 282298 561922 282366 561978
rect 282422 561922 312714 561978
rect 312770 561922 312838 561978
rect 312894 561922 312962 561978
rect 313018 561922 313086 561978
rect 313142 561922 343434 561978
rect 343490 561922 343558 561978
rect 343614 561922 343682 561978
rect 343738 561922 343806 561978
rect 343862 561922 374154 561978
rect 374210 561922 374278 561978
rect 374334 561922 374402 561978
rect 374458 561922 374526 561978
rect 374582 561922 404874 561978
rect 404930 561922 404998 561978
rect 405054 561922 405122 561978
rect 405178 561922 405246 561978
rect 405302 561922 435594 561978
rect 435650 561922 435718 561978
rect 435774 561922 435842 561978
rect 435898 561922 435966 561978
rect 436022 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect 4156 557938 459524 557954
rect 4156 557882 4172 557938
rect 4228 557882 459452 557938
rect 459508 557882 459524 557938
rect 4156 557866 459524 557882
rect 4156 551278 452804 551294
rect 4156 551222 4172 551278
rect 4228 551222 452732 551278
rect 452788 551222 452804 551278
rect 4156 551206 452804 551222
rect 55340 551098 590676 551114
rect 55340 551042 55356 551098
rect 55412 551042 590604 551098
rect 590660 551042 590676 551098
rect 55340 551026 590676 551042
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 179878 550350
rect 179934 550294 180002 550350
rect 180058 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 210598 550350
rect 210654 550294 210722 550350
rect 210778 550294 224274 550350
rect 224330 550294 224398 550350
rect 224454 550294 224522 550350
rect 224578 550294 224646 550350
rect 224702 550294 254994 550350
rect 255050 550294 255118 550350
rect 255174 550294 255242 550350
rect 255298 550294 255366 550350
rect 255422 550294 285714 550350
rect 285770 550294 285838 550350
rect 285894 550294 285962 550350
rect 286018 550294 286086 550350
rect 286142 550294 316434 550350
rect 316490 550294 316558 550350
rect 316614 550294 316682 550350
rect 316738 550294 316806 550350
rect 316862 550294 347154 550350
rect 347210 550294 347278 550350
rect 347334 550294 347402 550350
rect 347458 550294 347526 550350
rect 347582 550294 377874 550350
rect 377930 550294 377998 550350
rect 378054 550294 378122 550350
rect 378178 550294 378246 550350
rect 378302 550294 408594 550350
rect 408650 550294 408718 550350
rect 408774 550294 408842 550350
rect 408898 550294 408966 550350
rect 409022 550294 439314 550350
rect 439370 550294 439438 550350
rect 439494 550294 439562 550350
rect 439618 550294 439686 550350
rect 439742 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 179878 550226
rect 179934 550170 180002 550226
rect 180058 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 210598 550226
rect 210654 550170 210722 550226
rect 210778 550170 224274 550226
rect 224330 550170 224398 550226
rect 224454 550170 224522 550226
rect 224578 550170 224646 550226
rect 224702 550170 254994 550226
rect 255050 550170 255118 550226
rect 255174 550170 255242 550226
rect 255298 550170 255366 550226
rect 255422 550170 285714 550226
rect 285770 550170 285838 550226
rect 285894 550170 285962 550226
rect 286018 550170 286086 550226
rect 286142 550170 316434 550226
rect 316490 550170 316558 550226
rect 316614 550170 316682 550226
rect 316738 550170 316806 550226
rect 316862 550170 347154 550226
rect 347210 550170 347278 550226
rect 347334 550170 347402 550226
rect 347458 550170 347526 550226
rect 347582 550170 377874 550226
rect 377930 550170 377998 550226
rect 378054 550170 378122 550226
rect 378178 550170 378246 550226
rect 378302 550170 408594 550226
rect 408650 550170 408718 550226
rect 408774 550170 408842 550226
rect 408898 550170 408966 550226
rect 409022 550170 439314 550226
rect 439370 550170 439438 550226
rect 439494 550170 439562 550226
rect 439618 550170 439686 550226
rect 439742 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 179878 550102
rect 179934 550046 180002 550102
rect 180058 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 210598 550102
rect 210654 550046 210722 550102
rect 210778 550046 224274 550102
rect 224330 550046 224398 550102
rect 224454 550046 224522 550102
rect 224578 550046 224646 550102
rect 224702 550046 254994 550102
rect 255050 550046 255118 550102
rect 255174 550046 255242 550102
rect 255298 550046 255366 550102
rect 255422 550046 285714 550102
rect 285770 550046 285838 550102
rect 285894 550046 285962 550102
rect 286018 550046 286086 550102
rect 286142 550046 316434 550102
rect 316490 550046 316558 550102
rect 316614 550046 316682 550102
rect 316738 550046 316806 550102
rect 316862 550046 347154 550102
rect 347210 550046 347278 550102
rect 347334 550046 347402 550102
rect 347458 550046 347526 550102
rect 347582 550046 377874 550102
rect 377930 550046 377998 550102
rect 378054 550046 378122 550102
rect 378178 550046 378246 550102
rect 378302 550046 408594 550102
rect 408650 550046 408718 550102
rect 408774 550046 408842 550102
rect 408898 550046 408966 550102
rect 409022 550046 439314 550102
rect 439370 550046 439438 550102
rect 439494 550046 439562 550102
rect 439618 550046 439686 550102
rect 439742 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 179878 549978
rect 179934 549922 180002 549978
rect 180058 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 210598 549978
rect 210654 549922 210722 549978
rect 210778 549922 224274 549978
rect 224330 549922 224398 549978
rect 224454 549922 224522 549978
rect 224578 549922 224646 549978
rect 224702 549922 254994 549978
rect 255050 549922 255118 549978
rect 255174 549922 255242 549978
rect 255298 549922 255366 549978
rect 255422 549922 285714 549978
rect 285770 549922 285838 549978
rect 285894 549922 285962 549978
rect 286018 549922 286086 549978
rect 286142 549922 316434 549978
rect 316490 549922 316558 549978
rect 316614 549922 316682 549978
rect 316738 549922 316806 549978
rect 316862 549922 347154 549978
rect 347210 549922 347278 549978
rect 347334 549922 347402 549978
rect 347458 549922 347526 549978
rect 347582 549922 377874 549978
rect 377930 549922 377998 549978
rect 378054 549922 378122 549978
rect 378178 549922 378246 549978
rect 378302 549922 408594 549978
rect 408650 549922 408718 549978
rect 408774 549922 408842 549978
rect 408898 549922 408966 549978
rect 409022 549922 439314 549978
rect 439370 549922 439438 549978
rect 439494 549922 439562 549978
rect 439618 549922 439686 549978
rect 439742 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect 4268 548218 457844 548234
rect 4268 548162 4284 548218
rect 4340 548162 457772 548218
rect 457828 548162 457844 548218
rect 4268 548146 457844 548162
rect 121980 548038 590564 548054
rect 121980 547982 121996 548038
rect 122052 547982 590492 548038
rect 590548 547982 590564 548038
rect 121980 547966 590564 547982
rect 58700 547858 590228 547874
rect 58700 547802 58716 547858
rect 58772 547802 590156 547858
rect 590212 547802 590228 547858
rect 58700 547786 590228 547802
rect 268700 546418 556292 546434
rect 268700 546362 268716 546418
rect 268772 546362 556220 546418
rect 556276 546362 556292 546418
rect 268700 546346 556292 546362
rect 267020 546238 556180 546254
rect 267020 546182 267036 546238
rect 267092 546182 556108 546238
rect 556164 546182 556180 546238
rect 267020 546166 556180 546182
rect -1916 544433 597980 544446
rect -1916 544377 94810 544433
rect 94866 544377 94934 544433
rect 94990 544377 95058 544433
rect 95114 544377 95182 544433
rect 95238 544377 95306 544433
rect 95362 544377 95430 544433
rect 95486 544377 95554 544433
rect 95610 544377 95678 544433
rect 95734 544377 95802 544433
rect 95858 544377 95926 544433
rect 95982 544377 96050 544433
rect 96106 544377 96174 544433
rect 96230 544377 96298 544433
rect 96354 544377 96422 544433
rect 96478 544377 96546 544433
rect 96602 544377 96670 544433
rect 96726 544377 96794 544433
rect 96850 544377 96918 544433
rect 96974 544377 97042 544433
rect 97098 544377 97166 544433
rect 97222 544377 97290 544433
rect 97346 544377 97414 544433
rect 97470 544377 97538 544433
rect 97594 544377 97662 544433
rect 97718 544377 97786 544433
rect 97842 544377 97910 544433
rect 97966 544377 98034 544433
rect 98090 544377 98158 544433
rect 98214 544377 98282 544433
rect 98338 544377 98406 544433
rect 98462 544377 98530 544433
rect 98586 544377 98654 544433
rect 98710 544377 98778 544433
rect 98834 544377 98902 544433
rect 98958 544377 99026 544433
rect 99082 544377 99150 544433
rect 99206 544377 99274 544433
rect 99330 544377 99398 544433
rect 99454 544377 99522 544433
rect 99578 544377 99646 544433
rect 99702 544377 99770 544433
rect 99826 544377 99894 544433
rect 99950 544377 100018 544433
rect 100074 544377 100142 544433
rect 100198 544377 100266 544433
rect 100322 544377 100390 544433
rect 100446 544377 100514 544433
rect 100570 544377 100638 544433
rect 100694 544377 100762 544433
rect 100818 544377 100886 544433
rect 100942 544377 101010 544433
rect 101066 544377 101134 544433
rect 101190 544377 101258 544433
rect 101314 544377 101382 544433
rect 101438 544377 101506 544433
rect 101562 544377 101630 544433
rect 101686 544377 101754 544433
rect 101810 544377 101878 544433
rect 101934 544377 102002 544433
rect 102058 544377 102126 544433
rect 102182 544377 102250 544433
rect 102306 544377 102374 544433
rect 102430 544377 102498 544433
rect 102554 544377 102622 544433
rect 102678 544377 102746 544433
rect 102802 544377 102870 544433
rect 102926 544377 102994 544433
rect 103050 544377 103118 544433
rect 103174 544377 103242 544433
rect 103298 544377 103366 544433
rect 103422 544377 103490 544433
rect 103546 544377 103614 544433
rect 103670 544377 103738 544433
rect 103794 544377 103862 544433
rect 103918 544377 103986 544433
rect 104042 544377 104110 544433
rect 104166 544377 104234 544433
rect 104290 544377 104358 544433
rect 104414 544377 104482 544433
rect 104538 544377 104606 544433
rect 104662 544377 104730 544433
rect 104786 544377 104854 544433
rect 104910 544377 104978 544433
rect 105034 544377 105102 544433
rect 105158 544377 105226 544433
rect 105282 544377 105350 544433
rect 105406 544377 105474 544433
rect 105530 544377 105598 544433
rect 105654 544377 105722 544433
rect 105778 544377 105846 544433
rect 105902 544377 105970 544433
rect 106026 544377 106094 544433
rect 106150 544377 106218 544433
rect 106274 544377 106342 544433
rect 106398 544377 106466 544433
rect 106522 544377 106590 544433
rect 106646 544377 106714 544433
rect 106770 544377 106838 544433
rect 106894 544377 106962 544433
rect 107018 544377 107086 544433
rect 107142 544377 107210 544433
rect 107266 544377 107334 544433
rect 107390 544377 597980 544433
rect -1916 544350 597980 544377
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544309 128394 544350
rect 67382 544294 94810 544309
rect -1916 544253 94810 544294
rect 94866 544253 94934 544309
rect 94990 544253 95058 544309
rect 95114 544253 95182 544309
rect 95238 544253 95306 544309
rect 95362 544253 95430 544309
rect 95486 544253 95554 544309
rect 95610 544253 95678 544309
rect 95734 544253 95802 544309
rect 95858 544253 95926 544309
rect 95982 544253 96050 544309
rect 96106 544253 96174 544309
rect 96230 544253 96298 544309
rect 96354 544253 96422 544309
rect 96478 544253 96546 544309
rect 96602 544253 96670 544309
rect 96726 544253 96794 544309
rect 96850 544253 96918 544309
rect 96974 544253 97042 544309
rect 97098 544253 97166 544309
rect 97222 544253 97290 544309
rect 97346 544253 97414 544309
rect 97470 544253 97538 544309
rect 97594 544253 97662 544309
rect 97718 544253 97786 544309
rect 97842 544253 97910 544309
rect 97966 544253 98034 544309
rect 98090 544253 98158 544309
rect 98214 544253 98282 544309
rect 98338 544253 98406 544309
rect 98462 544253 98530 544309
rect 98586 544253 98654 544309
rect 98710 544253 98778 544309
rect 98834 544253 98902 544309
rect 98958 544253 99026 544309
rect 99082 544253 99150 544309
rect 99206 544253 99274 544309
rect 99330 544253 99398 544309
rect 99454 544253 99522 544309
rect 99578 544253 99646 544309
rect 99702 544253 99770 544309
rect 99826 544253 99894 544309
rect 99950 544253 100018 544309
rect 100074 544253 100142 544309
rect 100198 544253 100266 544309
rect 100322 544253 100390 544309
rect 100446 544253 100514 544309
rect 100570 544253 100638 544309
rect 100694 544253 100762 544309
rect 100818 544253 100886 544309
rect 100942 544253 101010 544309
rect 101066 544253 101134 544309
rect 101190 544253 101258 544309
rect 101314 544253 101382 544309
rect 101438 544253 101506 544309
rect 101562 544253 101630 544309
rect 101686 544253 101754 544309
rect 101810 544253 101878 544309
rect 101934 544253 102002 544309
rect 102058 544253 102126 544309
rect 102182 544253 102250 544309
rect 102306 544253 102374 544309
rect 102430 544253 102498 544309
rect 102554 544253 102622 544309
rect 102678 544253 102746 544309
rect 102802 544253 102870 544309
rect 102926 544253 102994 544309
rect 103050 544253 103118 544309
rect 103174 544253 103242 544309
rect 103298 544253 103366 544309
rect 103422 544253 103490 544309
rect 103546 544253 103614 544309
rect 103670 544253 103738 544309
rect 103794 544253 103862 544309
rect 103918 544253 103986 544309
rect 104042 544253 104110 544309
rect 104166 544253 104234 544309
rect 104290 544253 104358 544309
rect 104414 544253 104482 544309
rect 104538 544253 104606 544309
rect 104662 544253 104730 544309
rect 104786 544253 104854 544309
rect 104910 544253 104978 544309
rect 105034 544253 105102 544309
rect 105158 544253 105226 544309
rect 105282 544253 105350 544309
rect 105406 544253 105474 544309
rect 105530 544253 105598 544309
rect 105654 544253 105722 544309
rect 105778 544253 105846 544309
rect 105902 544253 105970 544309
rect 106026 544253 106094 544309
rect 106150 544253 106218 544309
rect 106274 544253 106342 544309
rect 106398 544253 106466 544309
rect 106522 544253 106590 544309
rect 106646 544253 106714 544309
rect 106770 544253 106838 544309
rect 106894 544253 106962 544309
rect 107018 544253 107086 544309
rect 107142 544253 107210 544309
rect 107266 544253 107334 544309
rect 107390 544294 128394 544309
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 164518 544350
rect 164574 544294 164642 544350
rect 164698 544294 195238 544350
rect 195294 544294 195362 544350
rect 195418 544294 220554 544350
rect 220610 544294 220678 544350
rect 220734 544294 220802 544350
rect 220858 544294 220926 544350
rect 220982 544294 251274 544350
rect 251330 544294 251398 544350
rect 251454 544294 251522 544350
rect 251578 544294 251646 544350
rect 251702 544294 281994 544350
rect 282050 544294 282118 544350
rect 282174 544294 282242 544350
rect 282298 544294 282366 544350
rect 282422 544294 304518 544350
rect 304574 544294 304642 544350
rect 304698 544294 335238 544350
rect 335294 544294 335362 544350
rect 335418 544294 365958 544350
rect 366014 544294 366082 544350
rect 366138 544294 396678 544350
rect 396734 544294 396802 544350
rect 396858 544294 427398 544350
rect 427454 544294 427522 544350
rect 427578 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect 107390 544253 597980 544294
rect -1916 544226 597980 544253
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 164518 544226
rect 164574 544170 164642 544226
rect 164698 544170 195238 544226
rect 195294 544170 195362 544226
rect 195418 544170 220554 544226
rect 220610 544170 220678 544226
rect 220734 544170 220802 544226
rect 220858 544170 220926 544226
rect 220982 544170 251274 544226
rect 251330 544170 251398 544226
rect 251454 544170 251522 544226
rect 251578 544170 251646 544226
rect 251702 544170 281994 544226
rect 282050 544170 282118 544226
rect 282174 544170 282242 544226
rect 282298 544170 282366 544226
rect 282422 544170 304518 544226
rect 304574 544170 304642 544226
rect 304698 544170 335238 544226
rect 335294 544170 335362 544226
rect 335418 544170 365958 544226
rect 366014 544170 366082 544226
rect 366138 544170 396678 544226
rect 396734 544170 396802 544226
rect 396858 544170 427398 544226
rect 427454 544170 427522 544226
rect 427578 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544090 128394 544102
rect 67382 544046 94630 544090
rect -1916 544034 94630 544046
rect 94686 544034 94754 544090
rect 94810 544034 94878 544090
rect 94934 544034 95002 544090
rect 95058 544034 95126 544090
rect 95182 544034 95250 544090
rect 95306 544034 95374 544090
rect 95430 544034 95498 544090
rect 95554 544034 95622 544090
rect 95678 544034 95746 544090
rect 95802 544034 95870 544090
rect 95926 544034 95994 544090
rect 96050 544034 96118 544090
rect 96174 544034 96242 544090
rect 96298 544034 96366 544090
rect 96422 544034 96490 544090
rect 96546 544034 96614 544090
rect 96670 544034 96738 544090
rect 96794 544034 96862 544090
rect 96918 544034 96986 544090
rect 97042 544034 97110 544090
rect 97166 544034 97234 544090
rect 97290 544034 97358 544090
rect 97414 544034 97482 544090
rect 97538 544034 97606 544090
rect 97662 544034 97730 544090
rect 97786 544034 97854 544090
rect 97910 544034 97978 544090
rect 98034 544034 98102 544090
rect 98158 544034 98226 544090
rect 98282 544034 98350 544090
rect 98406 544034 98474 544090
rect 98530 544034 98598 544090
rect 98654 544034 98722 544090
rect 98778 544034 98846 544090
rect 98902 544034 98970 544090
rect 99026 544034 99094 544090
rect 99150 544034 99218 544090
rect 99274 544034 99342 544090
rect 99398 544034 99466 544090
rect 99522 544034 99590 544090
rect 99646 544034 99714 544090
rect 99770 544034 99838 544090
rect 99894 544034 99962 544090
rect 100018 544034 100086 544090
rect 100142 544034 100210 544090
rect 100266 544034 100334 544090
rect 100390 544034 100458 544090
rect 100514 544034 100582 544090
rect 100638 544034 100706 544090
rect 100762 544034 100830 544090
rect 100886 544034 100954 544090
rect 101010 544034 101078 544090
rect 101134 544034 101202 544090
rect 101258 544034 101326 544090
rect 101382 544034 101450 544090
rect 101506 544034 101574 544090
rect 101630 544034 101698 544090
rect 101754 544034 101822 544090
rect 101878 544034 101946 544090
rect 102002 544034 102070 544090
rect 102126 544034 102194 544090
rect 102250 544034 102318 544090
rect 102374 544034 102442 544090
rect 102498 544034 102566 544090
rect 102622 544034 102690 544090
rect 102746 544034 102814 544090
rect 102870 544034 102938 544090
rect 102994 544034 103062 544090
rect 103118 544034 103186 544090
rect 103242 544034 103310 544090
rect 103366 544034 103434 544090
rect 103490 544034 103558 544090
rect 103614 544034 103682 544090
rect 103738 544034 103806 544090
rect 103862 544034 103930 544090
rect 103986 544034 104054 544090
rect 104110 544034 104178 544090
rect 104234 544034 104302 544090
rect 104358 544034 104426 544090
rect 104482 544034 104550 544090
rect 104606 544034 104674 544090
rect 104730 544034 104798 544090
rect 104854 544034 104922 544090
rect 104978 544034 105046 544090
rect 105102 544034 105170 544090
rect 105226 544034 105294 544090
rect 105350 544034 105418 544090
rect 105474 544034 105542 544090
rect 105598 544034 105666 544090
rect 105722 544034 105790 544090
rect 105846 544034 105914 544090
rect 105970 544034 106038 544090
rect 106094 544034 106162 544090
rect 106218 544034 106286 544090
rect 106342 544034 106410 544090
rect 106466 544034 106534 544090
rect 106590 544034 106658 544090
rect 106714 544034 106782 544090
rect 106838 544034 106906 544090
rect 106962 544034 107030 544090
rect 107086 544034 107154 544090
rect 107210 544046 128394 544090
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 164518 544102
rect 164574 544046 164642 544102
rect 164698 544046 195238 544102
rect 195294 544046 195362 544102
rect 195418 544046 220554 544102
rect 220610 544046 220678 544102
rect 220734 544046 220802 544102
rect 220858 544046 220926 544102
rect 220982 544046 251274 544102
rect 251330 544046 251398 544102
rect 251454 544046 251522 544102
rect 251578 544046 251646 544102
rect 251702 544046 281994 544102
rect 282050 544046 282118 544102
rect 282174 544046 282242 544102
rect 282298 544046 282366 544102
rect 282422 544046 304518 544102
rect 304574 544046 304642 544102
rect 304698 544046 335238 544102
rect 335294 544046 335362 544102
rect 335418 544046 365958 544102
rect 366014 544046 366082 544102
rect 366138 544046 396678 544102
rect 396734 544046 396802 544102
rect 396858 544046 427398 544102
rect 427454 544046 427522 544102
rect 427578 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect 107210 544034 597980 544046
rect -1916 543978 597980 544034
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543966 128394 543978
rect 67382 543922 94630 543966
rect -1916 543910 94630 543922
rect 94686 543910 94754 543966
rect 94810 543910 94878 543966
rect 94934 543910 95002 543966
rect 95058 543910 95126 543966
rect 95182 543910 95250 543966
rect 95306 543910 95374 543966
rect 95430 543910 95498 543966
rect 95554 543910 95622 543966
rect 95678 543910 95746 543966
rect 95802 543910 95870 543966
rect 95926 543910 95994 543966
rect 96050 543910 96118 543966
rect 96174 543910 96242 543966
rect 96298 543910 96366 543966
rect 96422 543910 96490 543966
rect 96546 543910 96614 543966
rect 96670 543910 96738 543966
rect 96794 543910 96862 543966
rect 96918 543910 96986 543966
rect 97042 543910 97110 543966
rect 97166 543910 97234 543966
rect 97290 543910 97358 543966
rect 97414 543910 97482 543966
rect 97538 543910 97606 543966
rect 97662 543910 97730 543966
rect 97786 543910 97854 543966
rect 97910 543910 97978 543966
rect 98034 543910 98102 543966
rect 98158 543910 98226 543966
rect 98282 543910 98350 543966
rect 98406 543910 98474 543966
rect 98530 543910 98598 543966
rect 98654 543910 98722 543966
rect 98778 543910 98846 543966
rect 98902 543910 98970 543966
rect 99026 543910 99094 543966
rect 99150 543910 99218 543966
rect 99274 543910 99342 543966
rect 99398 543910 99466 543966
rect 99522 543910 99590 543966
rect 99646 543910 99714 543966
rect 99770 543910 99838 543966
rect 99894 543910 99962 543966
rect 100018 543910 100086 543966
rect 100142 543910 100210 543966
rect 100266 543910 100334 543966
rect 100390 543910 100458 543966
rect 100514 543910 100582 543966
rect 100638 543910 100706 543966
rect 100762 543910 100830 543966
rect 100886 543910 100954 543966
rect 101010 543910 101078 543966
rect 101134 543910 101202 543966
rect 101258 543910 101326 543966
rect 101382 543910 101450 543966
rect 101506 543910 101574 543966
rect 101630 543910 101698 543966
rect 101754 543910 101822 543966
rect 101878 543910 101946 543966
rect 102002 543910 102070 543966
rect 102126 543910 102194 543966
rect 102250 543910 102318 543966
rect 102374 543910 102442 543966
rect 102498 543910 102566 543966
rect 102622 543910 102690 543966
rect 102746 543910 102814 543966
rect 102870 543910 102938 543966
rect 102994 543910 103062 543966
rect 103118 543910 103186 543966
rect 103242 543910 103310 543966
rect 103366 543910 103434 543966
rect 103490 543910 103558 543966
rect 103614 543910 103682 543966
rect 103738 543910 103806 543966
rect 103862 543910 103930 543966
rect 103986 543910 104054 543966
rect 104110 543910 104178 543966
rect 104234 543910 104302 543966
rect 104358 543910 104426 543966
rect 104482 543910 104550 543966
rect 104606 543910 104674 543966
rect 104730 543910 104798 543966
rect 104854 543910 104922 543966
rect 104978 543910 105046 543966
rect 105102 543910 105170 543966
rect 105226 543910 105294 543966
rect 105350 543910 105418 543966
rect 105474 543910 105542 543966
rect 105598 543910 105666 543966
rect 105722 543910 105790 543966
rect 105846 543910 105914 543966
rect 105970 543910 106038 543966
rect 106094 543910 106162 543966
rect 106218 543910 106286 543966
rect 106342 543910 106410 543966
rect 106466 543910 106534 543966
rect 106590 543910 106658 543966
rect 106714 543910 106782 543966
rect 106838 543910 106906 543966
rect 106962 543910 107030 543966
rect 107086 543910 107154 543966
rect 107210 543922 128394 543966
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 164518 543978
rect 164574 543922 164642 543978
rect 164698 543922 195238 543978
rect 195294 543922 195362 543978
rect 195418 543922 220554 543978
rect 220610 543922 220678 543978
rect 220734 543922 220802 543978
rect 220858 543922 220926 543978
rect 220982 543922 251274 543978
rect 251330 543922 251398 543978
rect 251454 543922 251522 543978
rect 251578 543922 251646 543978
rect 251702 543922 281994 543978
rect 282050 543922 282118 543978
rect 282174 543922 282242 543978
rect 282298 543922 282366 543978
rect 282422 543922 304518 543978
rect 304574 543922 304642 543978
rect 304698 543922 335238 543978
rect 335294 543922 335362 543978
rect 335418 543922 365958 543978
rect 366014 543922 366082 543978
rect 366138 543922 396678 543978
rect 396734 543922 396802 543978
rect 396858 543922 427398 543978
rect 427454 543922 427522 543978
rect 427578 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect 107210 543910 597980 543922
rect -1916 543826 597980 543910
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532328 132114 532350
rect 40382 532294 68074 532328
rect -1916 532272 68074 532294
rect 68130 532272 68198 532328
rect 68254 532272 68322 532328
rect 68378 532272 68446 532328
rect 68502 532272 68570 532328
rect 68626 532272 68694 532328
rect 68750 532272 68818 532328
rect 68874 532272 68942 532328
rect 68998 532272 69066 532328
rect 69122 532272 69190 532328
rect 69246 532272 69314 532328
rect 69370 532272 69438 532328
rect 69494 532272 69562 532328
rect 69618 532272 69686 532328
rect 69742 532272 69810 532328
rect 69866 532272 69934 532328
rect 69990 532272 70058 532328
rect 70114 532272 70182 532328
rect 70238 532272 70306 532328
rect 70362 532272 70430 532328
rect 70486 532272 70554 532328
rect 70610 532272 70678 532328
rect 70734 532272 70802 532328
rect 70858 532272 70926 532328
rect 70982 532272 71050 532328
rect 71106 532272 71174 532328
rect 71230 532272 71298 532328
rect 71354 532272 71422 532328
rect 71478 532272 71546 532328
rect 71602 532272 71670 532328
rect 71726 532272 71794 532328
rect 71850 532272 71918 532328
rect 71974 532272 72042 532328
rect 72098 532272 72166 532328
rect 72222 532272 72290 532328
rect 72346 532272 72414 532328
rect 72470 532272 72538 532328
rect 72594 532272 72662 532328
rect 72718 532272 72786 532328
rect 72842 532272 72910 532328
rect 72966 532272 73034 532328
rect 73090 532272 73158 532328
rect 73214 532272 73282 532328
rect 73338 532272 73406 532328
rect 73462 532272 73530 532328
rect 73586 532272 73654 532328
rect 73710 532272 73778 532328
rect 73834 532272 73902 532328
rect 73958 532272 74026 532328
rect 74082 532272 74150 532328
rect 74206 532272 74274 532328
rect 74330 532272 74398 532328
rect 74454 532272 74522 532328
rect 74578 532272 74646 532328
rect 74702 532272 74770 532328
rect 74826 532272 74894 532328
rect 74950 532272 75018 532328
rect 75074 532272 75142 532328
rect 75198 532272 75266 532328
rect 75322 532272 75390 532328
rect 75446 532294 132114 532328
rect 132170 532294 132238 532350
rect 132294 532294 132362 532350
rect 132418 532294 132486 532350
rect 132542 532294 179878 532350
rect 179934 532294 180002 532350
rect 180058 532294 210598 532350
rect 210654 532294 210722 532350
rect 210778 532294 224274 532350
rect 224330 532294 224398 532350
rect 224454 532294 224522 532350
rect 224578 532294 224646 532350
rect 224702 532294 254994 532350
rect 255050 532294 255118 532350
rect 255174 532294 255242 532350
rect 255298 532294 255366 532350
rect 255422 532294 285714 532350
rect 285770 532294 285838 532350
rect 285894 532294 285962 532350
rect 286018 532294 286086 532350
rect 286142 532294 319878 532350
rect 319934 532294 320002 532350
rect 320058 532294 350598 532350
rect 350654 532294 350722 532350
rect 350778 532294 381318 532350
rect 381374 532294 381442 532350
rect 381498 532294 412038 532350
rect 412094 532294 412162 532350
rect 412218 532294 442758 532350
rect 442814 532294 442882 532350
rect 442938 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 75446 532272 597980 532294
rect -1916 532226 597980 532272
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 132114 532226
rect 132170 532170 132238 532226
rect 132294 532170 132362 532226
rect 132418 532170 132486 532226
rect 132542 532170 179878 532226
rect 179934 532170 180002 532226
rect 180058 532170 210598 532226
rect 210654 532170 210722 532226
rect 210778 532170 224274 532226
rect 224330 532170 224398 532226
rect 224454 532170 224522 532226
rect 224578 532170 224646 532226
rect 224702 532170 254994 532226
rect 255050 532170 255118 532226
rect 255174 532170 255242 532226
rect 255298 532170 255366 532226
rect 255422 532170 285714 532226
rect 285770 532170 285838 532226
rect 285894 532170 285962 532226
rect 286018 532170 286086 532226
rect 286142 532170 319878 532226
rect 319934 532170 320002 532226
rect 320058 532170 350598 532226
rect 350654 532170 350722 532226
rect 350778 532170 381318 532226
rect 381374 532170 381442 532226
rect 381498 532170 412038 532226
rect 412094 532170 412162 532226
rect 412218 532170 442758 532226
rect 442814 532170 442882 532226
rect 442938 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 132114 532102
rect 132170 532046 132238 532102
rect 132294 532046 132362 532102
rect 132418 532046 132486 532102
rect 132542 532046 179878 532102
rect 179934 532046 180002 532102
rect 180058 532046 210598 532102
rect 210654 532046 210722 532102
rect 210778 532046 224274 532102
rect 224330 532046 224398 532102
rect 224454 532046 224522 532102
rect 224578 532046 224646 532102
rect 224702 532046 254994 532102
rect 255050 532046 255118 532102
rect 255174 532046 255242 532102
rect 255298 532046 255366 532102
rect 255422 532046 285714 532102
rect 285770 532046 285838 532102
rect 285894 532046 285962 532102
rect 286018 532046 286086 532102
rect 286142 532046 319878 532102
rect 319934 532046 320002 532102
rect 320058 532046 350598 532102
rect 350654 532046 350722 532102
rect 350778 532046 381318 532102
rect 381374 532046 381442 532102
rect 381498 532046 412038 532102
rect 412094 532046 412162 532102
rect 412218 532046 442758 532102
rect 442814 532046 442882 532102
rect 442938 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 132114 531978
rect 132170 531922 132238 531978
rect 132294 531922 132362 531978
rect 132418 531922 132486 531978
rect 132542 531922 179878 531978
rect 179934 531922 180002 531978
rect 180058 531922 210598 531978
rect 210654 531922 210722 531978
rect 210778 531922 224274 531978
rect 224330 531922 224398 531978
rect 224454 531922 224522 531978
rect 224578 531922 224646 531978
rect 224702 531922 254994 531978
rect 255050 531922 255118 531978
rect 255174 531922 255242 531978
rect 255298 531922 255366 531978
rect 255422 531922 285714 531978
rect 285770 531922 285838 531978
rect 285894 531922 285962 531978
rect 286018 531922 286086 531978
rect 286142 531922 319878 531978
rect 319934 531922 320002 531978
rect 320058 531922 350598 531978
rect 350654 531922 350722 531978
rect 350778 531922 381318 531978
rect 381374 531922 381442 531978
rect 381498 531922 412038 531978
rect 412094 531922 412162 531978
rect 412218 531922 442758 531978
rect 442814 531922 442882 531978
rect 442938 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526432 597980 526446
rect -1916 526376 497034 526432
rect 497090 526376 497158 526432
rect 497214 526376 497282 526432
rect 497338 526376 497406 526432
rect 497462 526376 527754 526432
rect 527810 526376 527878 526432
rect 527934 526376 528002 526432
rect 528058 526376 528126 526432
rect 528182 526376 597980 526432
rect -1916 526350 597980 526376
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526328 128394 526350
rect 36662 526294 84890 526328
rect -1916 526272 84890 526294
rect 84946 526272 85014 526328
rect 85070 526272 85138 526328
rect 85194 526272 85262 526328
rect 85318 526272 85386 526328
rect 85442 526272 85510 526328
rect 85566 526272 85634 526328
rect 85690 526272 85758 526328
rect 85814 526272 85882 526328
rect 85938 526272 86006 526328
rect 86062 526272 86130 526328
rect 86186 526272 86254 526328
rect 86310 526272 86378 526328
rect 86434 526272 86502 526328
rect 86558 526272 86626 526328
rect 86682 526272 86750 526328
rect 86806 526272 86874 526328
rect 86930 526272 86998 526328
rect 87054 526272 87122 526328
rect 87178 526272 87246 526328
rect 87302 526272 87370 526328
rect 87426 526272 87494 526328
rect 87550 526272 87618 526328
rect 87674 526272 87742 526328
rect 87798 526272 87866 526328
rect 87922 526272 87990 526328
rect 88046 526272 88114 526328
rect 88170 526272 88238 526328
rect 88294 526272 88362 526328
rect 88418 526272 88486 526328
rect 88542 526272 88610 526328
rect 88666 526272 88734 526328
rect 88790 526272 88858 526328
rect 88914 526272 88982 526328
rect 89038 526272 89106 526328
rect 89162 526272 89230 526328
rect 89286 526272 89354 526328
rect 89410 526272 89478 526328
rect 89534 526272 89602 526328
rect 89658 526272 89726 526328
rect 89782 526272 89850 526328
rect 89906 526272 89974 526328
rect 90030 526272 90098 526328
rect 90154 526272 90222 526328
rect 90278 526272 90346 526328
rect 90402 526272 90470 526328
rect 90526 526272 90594 526328
rect 90650 526272 90718 526328
rect 90774 526272 90842 526328
rect 90898 526272 90966 526328
rect 91022 526272 91090 526328
rect 91146 526272 91214 526328
rect 91270 526272 91338 526328
rect 91394 526272 91462 526328
rect 91518 526272 91586 526328
rect 91642 526272 91710 526328
rect 91766 526272 91834 526328
rect 91890 526272 91958 526328
rect 92014 526272 92082 526328
rect 92138 526272 92206 526328
rect 92262 526272 92330 526328
rect 92386 526272 92454 526328
rect 92510 526272 92578 526328
rect 92634 526272 92702 526328
rect 92758 526272 92826 526328
rect 92882 526272 92950 526328
rect 93006 526272 93074 526328
rect 93130 526272 93198 526328
rect 93254 526272 93322 526328
rect 93378 526272 93446 526328
rect 93502 526272 93570 526328
rect 93626 526272 93694 526328
rect 93750 526272 93818 526328
rect 93874 526272 93942 526328
rect 93998 526272 94066 526328
rect 94122 526272 94190 526328
rect 94246 526272 94314 526328
rect 94370 526272 94438 526328
rect 94494 526272 94562 526328
rect 94618 526272 94686 526328
rect 94742 526272 94810 526328
rect 94866 526272 94934 526328
rect 94990 526272 95058 526328
rect 95114 526272 95182 526328
rect 95238 526272 95306 526328
rect 95362 526272 95430 526328
rect 95486 526272 95554 526328
rect 95610 526272 95678 526328
rect 95734 526272 95802 526328
rect 95858 526272 95926 526328
rect 95982 526272 96050 526328
rect 96106 526272 96174 526328
rect 96230 526272 96298 526328
rect 96354 526272 96422 526328
rect 96478 526272 96546 526328
rect 96602 526272 96670 526328
rect 96726 526272 96794 526328
rect 96850 526272 96918 526328
rect 96974 526272 97042 526328
rect 97098 526272 97166 526328
rect 97222 526272 97290 526328
rect 97346 526272 97414 526328
rect 97470 526272 97538 526328
rect 97594 526272 97662 526328
rect 97718 526272 97786 526328
rect 97842 526272 97910 526328
rect 97966 526272 98034 526328
rect 98090 526272 98158 526328
rect 98214 526272 98282 526328
rect 98338 526272 98406 526328
rect 98462 526272 98530 526328
rect 98586 526272 98654 526328
rect 98710 526294 128394 526328
rect 128450 526294 128518 526350
rect 128574 526294 128642 526350
rect 128698 526294 128766 526350
rect 128822 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 164518 526350
rect 164574 526294 164642 526350
rect 164698 526294 195238 526350
rect 195294 526294 195362 526350
rect 195418 526294 220554 526350
rect 220610 526294 220678 526350
rect 220734 526294 220802 526350
rect 220858 526294 220926 526350
rect 220982 526294 251274 526350
rect 251330 526294 251398 526350
rect 251454 526294 251522 526350
rect 251578 526294 251646 526350
rect 251702 526294 281994 526350
rect 282050 526294 282118 526350
rect 282174 526294 282242 526350
rect 282298 526294 282366 526350
rect 282422 526294 304518 526350
rect 304574 526294 304642 526350
rect 304698 526294 335238 526350
rect 335294 526294 335362 526350
rect 335418 526294 365958 526350
rect 366014 526294 366082 526350
rect 366138 526294 396678 526350
rect 396734 526294 396802 526350
rect 396858 526294 427398 526350
rect 427454 526294 427522 526350
rect 427578 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 474518 526350
rect 474574 526294 474642 526350
rect 474698 526308 505238 526350
rect 474698 526294 497034 526308
rect 98710 526272 497034 526294
rect -1916 526252 497034 526272
rect 497090 526252 497158 526308
rect 497214 526252 497282 526308
rect 497338 526252 497406 526308
rect 497462 526294 505238 526308
rect 505294 526294 505362 526350
rect 505418 526308 535958 526350
rect 505418 526294 527754 526308
rect 497462 526252 527754 526294
rect 527810 526252 527878 526308
rect 527934 526252 528002 526308
rect 528058 526252 528126 526308
rect 528182 526294 535958 526308
rect 536014 526294 536082 526350
rect 536138 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect 528182 526252 597980 526294
rect -1916 526226 597980 526252
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 128394 526226
rect 128450 526170 128518 526226
rect 128574 526170 128642 526226
rect 128698 526170 128766 526226
rect 128822 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 164518 526226
rect 164574 526170 164642 526226
rect 164698 526170 195238 526226
rect 195294 526170 195362 526226
rect 195418 526170 220554 526226
rect 220610 526170 220678 526226
rect 220734 526170 220802 526226
rect 220858 526170 220926 526226
rect 220982 526170 251274 526226
rect 251330 526170 251398 526226
rect 251454 526170 251522 526226
rect 251578 526170 251646 526226
rect 251702 526170 281994 526226
rect 282050 526170 282118 526226
rect 282174 526170 282242 526226
rect 282298 526170 282366 526226
rect 282422 526170 304518 526226
rect 304574 526170 304642 526226
rect 304698 526170 335238 526226
rect 335294 526170 335362 526226
rect 335418 526170 365958 526226
rect 366014 526170 366082 526226
rect 366138 526170 396678 526226
rect 396734 526170 396802 526226
rect 396858 526170 427398 526226
rect 427454 526170 427522 526226
rect 427578 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 474518 526226
rect 474574 526170 474642 526226
rect 474698 526170 505238 526226
rect 505294 526170 505362 526226
rect 505418 526170 535958 526226
rect 536014 526170 536082 526226
rect 536138 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526090 128394 526102
rect 36662 526046 84772 526090
rect -1916 526034 84772 526046
rect 84828 526034 84896 526090
rect 84952 526034 85020 526090
rect 85076 526034 85144 526090
rect 85200 526034 85268 526090
rect 85324 526034 85392 526090
rect 85448 526034 85516 526090
rect 85572 526034 85640 526090
rect 85696 526034 85764 526090
rect 85820 526034 85888 526090
rect 85944 526034 86012 526090
rect 86068 526034 86136 526090
rect 86192 526034 86260 526090
rect 86316 526034 86384 526090
rect 86440 526034 86508 526090
rect 86564 526034 86632 526090
rect 86688 526034 86756 526090
rect 86812 526034 86880 526090
rect 86936 526034 87004 526090
rect 87060 526034 87128 526090
rect 87184 526034 87252 526090
rect 87308 526034 87376 526090
rect 87432 526034 87500 526090
rect 87556 526034 87624 526090
rect 87680 526034 87748 526090
rect 87804 526034 87872 526090
rect 87928 526034 87996 526090
rect 88052 526034 88120 526090
rect 88176 526034 88244 526090
rect 88300 526034 88368 526090
rect 88424 526034 88492 526090
rect 88548 526034 88616 526090
rect 88672 526034 88740 526090
rect 88796 526034 88864 526090
rect 88920 526034 88988 526090
rect 89044 526034 89112 526090
rect 89168 526034 89236 526090
rect 89292 526034 89360 526090
rect 89416 526034 89484 526090
rect 89540 526034 89608 526090
rect 89664 526034 89732 526090
rect 89788 526034 89856 526090
rect 89912 526034 89980 526090
rect 90036 526034 90104 526090
rect 90160 526034 90228 526090
rect 90284 526034 90352 526090
rect 90408 526034 90476 526090
rect 90532 526034 90600 526090
rect 90656 526034 90724 526090
rect 90780 526034 90848 526090
rect 90904 526034 90972 526090
rect 91028 526034 91096 526090
rect 91152 526034 91220 526090
rect 91276 526034 91344 526090
rect 91400 526034 91468 526090
rect 91524 526034 91592 526090
rect 91648 526034 91716 526090
rect 91772 526034 91840 526090
rect 91896 526034 91964 526090
rect 92020 526034 92088 526090
rect 92144 526034 92212 526090
rect 92268 526034 92336 526090
rect 92392 526034 92460 526090
rect 92516 526034 92584 526090
rect 92640 526034 92708 526090
rect 92764 526034 92832 526090
rect 92888 526034 92956 526090
rect 93012 526034 93080 526090
rect 93136 526034 93204 526090
rect 93260 526034 93328 526090
rect 93384 526034 93452 526090
rect 93508 526034 93576 526090
rect 93632 526034 93700 526090
rect 93756 526034 93824 526090
rect 93880 526034 93948 526090
rect 94004 526034 94072 526090
rect 94128 526034 94196 526090
rect 94252 526034 94320 526090
rect 94376 526034 94444 526090
rect 94500 526034 94568 526090
rect 94624 526034 94692 526090
rect 94748 526034 94816 526090
rect 94872 526034 94940 526090
rect 94996 526034 95064 526090
rect 95120 526034 95188 526090
rect 95244 526034 95312 526090
rect 95368 526034 95436 526090
rect 95492 526034 95560 526090
rect 95616 526034 95684 526090
rect 95740 526034 95808 526090
rect 95864 526034 95932 526090
rect 95988 526034 96056 526090
rect 96112 526034 96180 526090
rect 96236 526034 96304 526090
rect 96360 526034 96428 526090
rect 96484 526034 96552 526090
rect 96608 526034 96676 526090
rect 96732 526034 96800 526090
rect 96856 526034 96924 526090
rect 96980 526034 97048 526090
rect 97104 526034 97172 526090
rect 97228 526034 97296 526090
rect 97352 526034 97420 526090
rect 97476 526034 97544 526090
rect 97600 526034 97668 526090
rect 97724 526034 97792 526090
rect 97848 526034 97916 526090
rect 97972 526034 98040 526090
rect 98096 526034 98164 526090
rect 98220 526034 98288 526090
rect 98344 526034 98412 526090
rect 98468 526046 128394 526090
rect 128450 526046 128518 526102
rect 128574 526046 128642 526102
rect 128698 526046 128766 526102
rect 128822 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 164518 526102
rect 164574 526046 164642 526102
rect 164698 526046 195238 526102
rect 195294 526046 195362 526102
rect 195418 526046 220554 526102
rect 220610 526046 220678 526102
rect 220734 526046 220802 526102
rect 220858 526046 220926 526102
rect 220982 526046 251274 526102
rect 251330 526046 251398 526102
rect 251454 526046 251522 526102
rect 251578 526046 251646 526102
rect 251702 526046 281994 526102
rect 282050 526046 282118 526102
rect 282174 526046 282242 526102
rect 282298 526046 282366 526102
rect 282422 526046 304518 526102
rect 304574 526046 304642 526102
rect 304698 526046 335238 526102
rect 335294 526046 335362 526102
rect 335418 526046 365958 526102
rect 366014 526046 366082 526102
rect 366138 526046 396678 526102
rect 396734 526046 396802 526102
rect 396858 526046 427398 526102
rect 427454 526046 427522 526102
rect 427578 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 474518 526102
rect 474574 526046 474642 526102
rect 474698 526046 505238 526102
rect 505294 526046 505362 526102
rect 505418 526046 535958 526102
rect 536014 526046 536082 526102
rect 536138 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect 98468 526034 597980 526046
rect -1916 525978 597980 526034
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525966 128394 525978
rect 36662 525922 84772 525966
rect -1916 525910 84772 525922
rect 84828 525910 84896 525966
rect 84952 525910 85020 525966
rect 85076 525910 85144 525966
rect 85200 525910 85268 525966
rect 85324 525910 85392 525966
rect 85448 525910 85516 525966
rect 85572 525910 85640 525966
rect 85696 525910 85764 525966
rect 85820 525910 85888 525966
rect 85944 525910 86012 525966
rect 86068 525910 86136 525966
rect 86192 525910 86260 525966
rect 86316 525910 86384 525966
rect 86440 525910 86508 525966
rect 86564 525910 86632 525966
rect 86688 525910 86756 525966
rect 86812 525910 86880 525966
rect 86936 525910 87004 525966
rect 87060 525910 87128 525966
rect 87184 525910 87252 525966
rect 87308 525910 87376 525966
rect 87432 525910 87500 525966
rect 87556 525910 87624 525966
rect 87680 525910 87748 525966
rect 87804 525910 87872 525966
rect 87928 525910 87996 525966
rect 88052 525910 88120 525966
rect 88176 525910 88244 525966
rect 88300 525910 88368 525966
rect 88424 525910 88492 525966
rect 88548 525910 88616 525966
rect 88672 525910 88740 525966
rect 88796 525910 88864 525966
rect 88920 525910 88988 525966
rect 89044 525910 89112 525966
rect 89168 525910 89236 525966
rect 89292 525910 89360 525966
rect 89416 525910 89484 525966
rect 89540 525910 89608 525966
rect 89664 525910 89732 525966
rect 89788 525910 89856 525966
rect 89912 525910 89980 525966
rect 90036 525910 90104 525966
rect 90160 525910 90228 525966
rect 90284 525910 90352 525966
rect 90408 525910 90476 525966
rect 90532 525910 90600 525966
rect 90656 525910 90724 525966
rect 90780 525910 90848 525966
rect 90904 525910 90972 525966
rect 91028 525910 91096 525966
rect 91152 525910 91220 525966
rect 91276 525910 91344 525966
rect 91400 525910 91468 525966
rect 91524 525910 91592 525966
rect 91648 525910 91716 525966
rect 91772 525910 91840 525966
rect 91896 525910 91964 525966
rect 92020 525910 92088 525966
rect 92144 525910 92212 525966
rect 92268 525910 92336 525966
rect 92392 525910 92460 525966
rect 92516 525910 92584 525966
rect 92640 525910 92708 525966
rect 92764 525910 92832 525966
rect 92888 525910 92956 525966
rect 93012 525910 93080 525966
rect 93136 525910 93204 525966
rect 93260 525910 93328 525966
rect 93384 525910 93452 525966
rect 93508 525910 93576 525966
rect 93632 525910 93700 525966
rect 93756 525910 93824 525966
rect 93880 525910 93948 525966
rect 94004 525910 94072 525966
rect 94128 525910 94196 525966
rect 94252 525910 94320 525966
rect 94376 525910 94444 525966
rect 94500 525910 94568 525966
rect 94624 525910 94692 525966
rect 94748 525910 94816 525966
rect 94872 525910 94940 525966
rect 94996 525910 95064 525966
rect 95120 525910 95188 525966
rect 95244 525910 95312 525966
rect 95368 525910 95436 525966
rect 95492 525910 95560 525966
rect 95616 525910 95684 525966
rect 95740 525910 95808 525966
rect 95864 525910 95932 525966
rect 95988 525910 96056 525966
rect 96112 525910 96180 525966
rect 96236 525910 96304 525966
rect 96360 525910 96428 525966
rect 96484 525910 96552 525966
rect 96608 525910 96676 525966
rect 96732 525910 96800 525966
rect 96856 525910 96924 525966
rect 96980 525910 97048 525966
rect 97104 525910 97172 525966
rect 97228 525910 97296 525966
rect 97352 525910 97420 525966
rect 97476 525910 97544 525966
rect 97600 525910 97668 525966
rect 97724 525910 97792 525966
rect 97848 525910 97916 525966
rect 97972 525910 98040 525966
rect 98096 525910 98164 525966
rect 98220 525910 98288 525966
rect 98344 525910 98412 525966
rect 98468 525922 128394 525966
rect 128450 525922 128518 525978
rect 128574 525922 128642 525978
rect 128698 525922 128766 525978
rect 128822 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 164518 525978
rect 164574 525922 164642 525978
rect 164698 525922 195238 525978
rect 195294 525922 195362 525978
rect 195418 525922 220554 525978
rect 220610 525922 220678 525978
rect 220734 525922 220802 525978
rect 220858 525922 220926 525978
rect 220982 525922 251274 525978
rect 251330 525922 251398 525978
rect 251454 525922 251522 525978
rect 251578 525922 251646 525978
rect 251702 525922 281994 525978
rect 282050 525922 282118 525978
rect 282174 525922 282242 525978
rect 282298 525922 282366 525978
rect 282422 525922 304518 525978
rect 304574 525922 304642 525978
rect 304698 525922 335238 525978
rect 335294 525922 335362 525978
rect 335418 525922 365958 525978
rect 366014 525922 366082 525978
rect 366138 525922 396678 525978
rect 396734 525922 396802 525978
rect 396858 525922 427398 525978
rect 427454 525922 427522 525978
rect 427578 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 474518 525978
rect 474574 525922 474642 525978
rect 474698 525922 505238 525978
rect 505294 525922 505362 525978
rect 505418 525922 535958 525978
rect 536014 525922 536082 525978
rect 536138 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect 98468 525910 597980 525922
rect -1916 525826 597980 525910
rect 300508 521758 301940 521774
rect 300508 521702 300524 521758
rect 300580 521702 301868 521758
rect 301924 521702 301940 521758
rect 300508 521686 301940 521702
rect 300620 520318 301828 520334
rect 300620 520262 300636 520318
rect 300692 520262 301756 520318
rect 301812 520262 301828 520318
rect 300620 520246 301828 520262
rect 300508 516898 301716 516914
rect 300508 516842 300524 516898
rect 300580 516842 301644 516898
rect 301700 516842 301716 516898
rect 300508 516826 301716 516842
rect -1916 514412 597980 514446
rect -1916 514356 60026 514412
rect 60082 514356 60150 514412
rect 60206 514356 60274 514412
rect 60330 514356 60398 514412
rect 60454 514356 60522 514412
rect 60578 514356 60646 514412
rect 60702 514356 60770 514412
rect 60826 514356 60894 514412
rect 60950 514356 61018 514412
rect 61074 514356 61142 514412
rect 61198 514356 61266 514412
rect 61322 514356 61390 514412
rect 61446 514356 61514 514412
rect 61570 514356 61638 514412
rect 61694 514356 61762 514412
rect 61818 514356 61886 514412
rect 61942 514356 62010 514412
rect 62066 514356 62134 514412
rect 62190 514356 62258 514412
rect 62314 514356 62382 514412
rect 62438 514356 62506 514412
rect 62562 514356 62630 514412
rect 62686 514356 62754 514412
rect 62810 514356 62878 514412
rect 62934 514356 63002 514412
rect 63058 514356 63126 514412
rect 63182 514356 63250 514412
rect 63306 514356 63374 514412
rect 63430 514356 63498 514412
rect 63554 514356 63622 514412
rect 63678 514356 63746 514412
rect 63802 514356 63870 514412
rect 63926 514356 63994 514412
rect 64050 514356 64118 514412
rect 64174 514356 597980 514412
rect -1916 514350 597980 514356
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 132114 514350
rect 132170 514294 132238 514350
rect 132294 514294 132362 514350
rect 132418 514294 132486 514350
rect 132542 514294 179878 514350
rect 179934 514294 180002 514350
rect 180058 514294 210598 514350
rect 210654 514294 210722 514350
rect 210778 514294 224274 514350
rect 224330 514294 224398 514350
rect 224454 514294 224522 514350
rect 224578 514294 224646 514350
rect 224702 514294 254994 514350
rect 255050 514294 255118 514350
rect 255174 514294 255242 514350
rect 255298 514294 255366 514350
rect 255422 514294 285714 514350
rect 285770 514294 285838 514350
rect 285894 514294 285962 514350
rect 286018 514294 286086 514350
rect 286142 514294 319878 514350
rect 319934 514294 320002 514350
rect 320058 514294 350598 514350
rect 350654 514294 350722 514350
rect 350778 514294 381318 514350
rect 381374 514294 381442 514350
rect 381498 514294 412038 514350
rect 412094 514294 412162 514350
rect 412218 514294 442758 514350
rect 442814 514294 442882 514350
rect 442938 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 489878 514350
rect 489934 514294 490002 514350
rect 490058 514294 520598 514350
rect 520654 514294 520722 514350
rect 520778 514294 551318 514350
rect 551374 514294 551442 514350
rect 551498 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514288 597980 514294
rect -1916 514232 60026 514288
rect 60082 514232 60150 514288
rect 60206 514232 60274 514288
rect 60330 514232 60398 514288
rect 60454 514232 60522 514288
rect 60578 514232 60646 514288
rect 60702 514232 60770 514288
rect 60826 514232 60894 514288
rect 60950 514232 61018 514288
rect 61074 514232 61142 514288
rect 61198 514232 61266 514288
rect 61322 514232 61390 514288
rect 61446 514232 61514 514288
rect 61570 514232 61638 514288
rect 61694 514232 61762 514288
rect 61818 514232 61886 514288
rect 61942 514232 62010 514288
rect 62066 514232 62134 514288
rect 62190 514232 62258 514288
rect 62314 514232 62382 514288
rect 62438 514232 62506 514288
rect 62562 514232 62630 514288
rect 62686 514232 62754 514288
rect 62810 514232 62878 514288
rect 62934 514232 63002 514288
rect 63058 514232 63126 514288
rect 63182 514232 63250 514288
rect 63306 514232 63374 514288
rect 63430 514232 63498 514288
rect 63554 514232 63622 514288
rect 63678 514232 63746 514288
rect 63802 514232 63870 514288
rect 63926 514232 63994 514288
rect 64050 514232 64118 514288
rect 64174 514232 597980 514288
rect -1916 514226 597980 514232
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 132114 514226
rect 132170 514170 132238 514226
rect 132294 514170 132362 514226
rect 132418 514170 132486 514226
rect 132542 514170 179878 514226
rect 179934 514170 180002 514226
rect 180058 514170 210598 514226
rect 210654 514170 210722 514226
rect 210778 514170 224274 514226
rect 224330 514170 224398 514226
rect 224454 514170 224522 514226
rect 224578 514170 224646 514226
rect 224702 514170 254994 514226
rect 255050 514170 255118 514226
rect 255174 514170 255242 514226
rect 255298 514170 255366 514226
rect 255422 514170 285714 514226
rect 285770 514170 285838 514226
rect 285894 514170 285962 514226
rect 286018 514170 286086 514226
rect 286142 514170 319878 514226
rect 319934 514170 320002 514226
rect 320058 514170 350598 514226
rect 350654 514170 350722 514226
rect 350778 514170 381318 514226
rect 381374 514170 381442 514226
rect 381498 514170 412038 514226
rect 412094 514170 412162 514226
rect 412218 514170 442758 514226
rect 442814 514170 442882 514226
rect 442938 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 489878 514226
rect 489934 514170 490002 514226
rect 490058 514170 520598 514226
rect 520654 514170 520722 514226
rect 520778 514170 551318 514226
rect 551374 514170 551442 514226
rect 551498 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514164 597980 514170
rect -1916 514108 60026 514164
rect 60082 514108 60150 514164
rect 60206 514108 60274 514164
rect 60330 514108 60398 514164
rect 60454 514108 60522 514164
rect 60578 514108 60646 514164
rect 60702 514108 60770 514164
rect 60826 514108 60894 514164
rect 60950 514108 61018 514164
rect 61074 514108 61142 514164
rect 61198 514108 61266 514164
rect 61322 514108 61390 514164
rect 61446 514108 61514 514164
rect 61570 514108 61638 514164
rect 61694 514108 61762 514164
rect 61818 514108 61886 514164
rect 61942 514108 62010 514164
rect 62066 514108 62134 514164
rect 62190 514108 62258 514164
rect 62314 514108 62382 514164
rect 62438 514108 62506 514164
rect 62562 514108 62630 514164
rect 62686 514108 62754 514164
rect 62810 514108 62878 514164
rect 62934 514108 63002 514164
rect 63058 514108 63126 514164
rect 63182 514108 63250 514164
rect 63306 514108 63374 514164
rect 63430 514108 63498 514164
rect 63554 514108 63622 514164
rect 63678 514108 63746 514164
rect 63802 514108 63870 514164
rect 63926 514108 63994 514164
rect 64050 514108 64118 514164
rect 64174 514108 597980 514164
rect -1916 514102 597980 514108
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 132114 514102
rect 132170 514046 132238 514102
rect 132294 514046 132362 514102
rect 132418 514046 132486 514102
rect 132542 514046 179878 514102
rect 179934 514046 180002 514102
rect 180058 514046 210598 514102
rect 210654 514046 210722 514102
rect 210778 514046 224274 514102
rect 224330 514046 224398 514102
rect 224454 514046 224522 514102
rect 224578 514046 224646 514102
rect 224702 514046 254994 514102
rect 255050 514046 255118 514102
rect 255174 514046 255242 514102
rect 255298 514046 255366 514102
rect 255422 514046 285714 514102
rect 285770 514046 285838 514102
rect 285894 514046 285962 514102
rect 286018 514046 286086 514102
rect 286142 514046 319878 514102
rect 319934 514046 320002 514102
rect 320058 514046 350598 514102
rect 350654 514046 350722 514102
rect 350778 514046 381318 514102
rect 381374 514046 381442 514102
rect 381498 514046 412038 514102
rect 412094 514046 412162 514102
rect 412218 514046 442758 514102
rect 442814 514046 442882 514102
rect 442938 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 489878 514102
rect 489934 514046 490002 514102
rect 490058 514046 520598 514102
rect 520654 514046 520722 514102
rect 520778 514046 551318 514102
rect 551374 514046 551442 514102
rect 551498 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 514040 597980 514046
rect -1916 513984 60026 514040
rect 60082 513984 60150 514040
rect 60206 513984 60274 514040
rect 60330 513984 60398 514040
rect 60454 513984 60522 514040
rect 60578 513984 60646 514040
rect 60702 513984 60770 514040
rect 60826 513984 60894 514040
rect 60950 513984 61018 514040
rect 61074 513984 61142 514040
rect 61198 513984 61266 514040
rect 61322 513984 61390 514040
rect 61446 513984 61514 514040
rect 61570 513984 61638 514040
rect 61694 513984 61762 514040
rect 61818 513984 61886 514040
rect 61942 513984 62010 514040
rect 62066 513984 62134 514040
rect 62190 513984 62258 514040
rect 62314 513984 62382 514040
rect 62438 513984 62506 514040
rect 62562 513984 62630 514040
rect 62686 513984 62754 514040
rect 62810 513984 62878 514040
rect 62934 513984 63002 514040
rect 63058 513984 63126 514040
rect 63182 513984 63250 514040
rect 63306 513984 63374 514040
rect 63430 513984 63498 514040
rect 63554 513984 63622 514040
rect 63678 513984 63746 514040
rect 63802 513984 63870 514040
rect 63926 513984 63994 514040
rect 64050 513984 64118 514040
rect 64174 513984 597980 514040
rect -1916 513978 597980 513984
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 132114 513978
rect 132170 513922 132238 513978
rect 132294 513922 132362 513978
rect 132418 513922 132486 513978
rect 132542 513922 179878 513978
rect 179934 513922 180002 513978
rect 180058 513922 210598 513978
rect 210654 513922 210722 513978
rect 210778 513922 224274 513978
rect 224330 513922 224398 513978
rect 224454 513922 224522 513978
rect 224578 513922 224646 513978
rect 224702 513922 254994 513978
rect 255050 513922 255118 513978
rect 255174 513922 255242 513978
rect 255298 513922 255366 513978
rect 255422 513922 285714 513978
rect 285770 513922 285838 513978
rect 285894 513922 285962 513978
rect 286018 513922 286086 513978
rect 286142 513922 319878 513978
rect 319934 513922 320002 513978
rect 320058 513922 350598 513978
rect 350654 513922 350722 513978
rect 350778 513922 381318 513978
rect 381374 513922 381442 513978
rect 381498 513922 412038 513978
rect 412094 513922 412162 513978
rect 412218 513922 442758 513978
rect 442814 513922 442882 513978
rect 442938 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 489878 513978
rect 489934 513922 490002 513978
rect 490058 513922 520598 513978
rect 520654 513922 520722 513978
rect 520778 513922 551318 513978
rect 551374 513922 551442 513978
rect 551498 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513916 597980 513922
rect -1916 513860 60026 513916
rect 60082 513860 60150 513916
rect 60206 513860 60274 513916
rect 60330 513860 60398 513916
rect 60454 513860 60522 513916
rect 60578 513860 60646 513916
rect 60702 513860 60770 513916
rect 60826 513860 60894 513916
rect 60950 513860 61018 513916
rect 61074 513860 61142 513916
rect 61198 513860 61266 513916
rect 61322 513860 61390 513916
rect 61446 513860 61514 513916
rect 61570 513860 61638 513916
rect 61694 513860 61762 513916
rect 61818 513860 61886 513916
rect 61942 513860 62010 513916
rect 62066 513860 62134 513916
rect 62190 513860 62258 513916
rect 62314 513860 62382 513916
rect 62438 513860 62506 513916
rect 62562 513860 62630 513916
rect 62686 513860 62754 513916
rect 62810 513860 62878 513916
rect 62934 513860 63002 513916
rect 63058 513860 63126 513916
rect 63182 513860 63250 513916
rect 63306 513860 63374 513916
rect 63430 513860 63498 513916
rect 63554 513860 63622 513916
rect 63678 513860 63746 513916
rect 63802 513860 63870 513916
rect 63926 513860 63994 513916
rect 64050 513860 64118 513916
rect 64174 513860 597980 513916
rect -1916 513826 597980 513860
rect 300620 513658 301604 513674
rect 300620 513602 300636 513658
rect 300692 513602 301532 513658
rect 301588 513602 301604 513658
rect 300620 513586 301604 513602
rect -1916 508431 597980 508446
rect -1916 508375 78970 508431
rect 79026 508375 79094 508431
rect 79150 508375 79218 508431
rect 79274 508375 79342 508431
rect 79398 508375 79466 508431
rect 79522 508375 79590 508431
rect 79646 508375 79714 508431
rect 79770 508375 79838 508431
rect 79894 508375 79962 508431
rect 80018 508375 80086 508431
rect 80142 508375 80210 508431
rect 80266 508375 80334 508431
rect 80390 508375 80458 508431
rect 80514 508375 80582 508431
rect 80638 508375 80706 508431
rect 80762 508375 80830 508431
rect 80886 508375 80954 508431
rect 81010 508375 81078 508431
rect 81134 508375 81202 508431
rect 81258 508375 81326 508431
rect 81382 508375 81450 508431
rect 81506 508375 81574 508431
rect 81630 508375 81698 508431
rect 81754 508375 81822 508431
rect 81878 508375 81946 508431
rect 82002 508375 82070 508431
rect 82126 508375 82194 508431
rect 82250 508375 82318 508431
rect 82374 508375 82442 508431
rect 82498 508375 82566 508431
rect 82622 508375 82690 508431
rect 82746 508375 82814 508431
rect 82870 508375 82938 508431
rect 82994 508375 83062 508431
rect 83118 508375 83186 508431
rect 83242 508375 83310 508431
rect 83366 508375 83434 508431
rect 83490 508375 83558 508431
rect 83614 508375 83682 508431
rect 83738 508375 83806 508431
rect 83862 508375 83930 508431
rect 83986 508375 84054 508431
rect 84110 508375 597980 508431
rect -1916 508350 597980 508375
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 128394 508350
rect 128450 508294 128518 508350
rect 128574 508294 128642 508350
rect 128698 508294 128766 508350
rect 128822 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 164518 508350
rect 164574 508294 164642 508350
rect 164698 508294 195238 508350
rect 195294 508294 195362 508350
rect 195418 508294 220554 508350
rect 220610 508294 220678 508350
rect 220734 508294 220802 508350
rect 220858 508294 220926 508350
rect 220982 508294 251274 508350
rect 251330 508294 251398 508350
rect 251454 508294 251522 508350
rect 251578 508294 251646 508350
rect 251702 508294 281994 508350
rect 282050 508294 282118 508350
rect 282174 508294 282242 508350
rect 282298 508294 282366 508350
rect 282422 508294 304518 508350
rect 304574 508294 304642 508350
rect 304698 508294 335238 508350
rect 335294 508294 335362 508350
rect 335418 508294 365958 508350
rect 366014 508294 366082 508350
rect 366138 508294 396678 508350
rect 396734 508294 396802 508350
rect 396858 508294 427398 508350
rect 427454 508294 427522 508350
rect 427578 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 474518 508350
rect 474574 508294 474642 508350
rect 474698 508294 505238 508350
rect 505294 508294 505362 508350
rect 505418 508294 535958 508350
rect 536014 508294 536082 508350
rect 536138 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508208 128394 508226
rect 36662 508170 78850 508208
rect -1916 508152 78850 508170
rect 78906 508152 78974 508208
rect 79030 508152 79098 508208
rect 79154 508152 79222 508208
rect 79278 508152 79346 508208
rect 79402 508152 79470 508208
rect 79526 508152 79594 508208
rect 79650 508152 79718 508208
rect 79774 508152 79842 508208
rect 79898 508152 79966 508208
rect 80022 508152 80090 508208
rect 80146 508152 80214 508208
rect 80270 508152 80338 508208
rect 80394 508152 80462 508208
rect 80518 508152 80586 508208
rect 80642 508152 80710 508208
rect 80766 508152 80834 508208
rect 80890 508152 80958 508208
rect 81014 508152 81082 508208
rect 81138 508152 81206 508208
rect 81262 508152 81330 508208
rect 81386 508152 81454 508208
rect 81510 508152 81578 508208
rect 81634 508152 81702 508208
rect 81758 508152 81826 508208
rect 81882 508152 81950 508208
rect 82006 508152 82074 508208
rect 82130 508152 82198 508208
rect 82254 508152 82322 508208
rect 82378 508152 82446 508208
rect 82502 508152 82570 508208
rect 82626 508152 82694 508208
rect 82750 508152 82818 508208
rect 82874 508152 82942 508208
rect 82998 508152 83066 508208
rect 83122 508152 83190 508208
rect 83246 508152 83314 508208
rect 83370 508152 83438 508208
rect 83494 508152 83562 508208
rect 83618 508152 83686 508208
rect 83742 508152 83810 508208
rect 83866 508152 83934 508208
rect 83990 508170 128394 508208
rect 128450 508170 128518 508226
rect 128574 508170 128642 508226
rect 128698 508170 128766 508226
rect 128822 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 164518 508226
rect 164574 508170 164642 508226
rect 164698 508170 195238 508226
rect 195294 508170 195362 508226
rect 195418 508170 220554 508226
rect 220610 508170 220678 508226
rect 220734 508170 220802 508226
rect 220858 508170 220926 508226
rect 220982 508170 251274 508226
rect 251330 508170 251398 508226
rect 251454 508170 251522 508226
rect 251578 508170 251646 508226
rect 251702 508170 281994 508226
rect 282050 508170 282118 508226
rect 282174 508170 282242 508226
rect 282298 508170 282366 508226
rect 282422 508170 304518 508226
rect 304574 508170 304642 508226
rect 304698 508170 335238 508226
rect 335294 508170 335362 508226
rect 335418 508170 365958 508226
rect 366014 508170 366082 508226
rect 366138 508170 396678 508226
rect 396734 508170 396802 508226
rect 396858 508170 427398 508226
rect 427454 508170 427522 508226
rect 427578 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 474518 508226
rect 474574 508170 474642 508226
rect 474698 508170 505238 508226
rect 505294 508170 505362 508226
rect 505418 508170 535958 508226
rect 536014 508170 536082 508226
rect 536138 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect 83990 508152 597980 508170
rect -1916 508102 597980 508152
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 128394 508102
rect 128450 508046 128518 508102
rect 128574 508046 128642 508102
rect 128698 508046 128766 508102
rect 128822 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 164518 508102
rect 164574 508046 164642 508102
rect 164698 508046 195238 508102
rect 195294 508046 195362 508102
rect 195418 508046 220554 508102
rect 220610 508046 220678 508102
rect 220734 508046 220802 508102
rect 220858 508046 220926 508102
rect 220982 508046 251274 508102
rect 251330 508046 251398 508102
rect 251454 508046 251522 508102
rect 251578 508046 251646 508102
rect 251702 508046 281994 508102
rect 282050 508046 282118 508102
rect 282174 508046 282242 508102
rect 282298 508046 282366 508102
rect 282422 508046 304518 508102
rect 304574 508046 304642 508102
rect 304698 508046 335238 508102
rect 335294 508046 335362 508102
rect 335418 508046 365958 508102
rect 366014 508046 366082 508102
rect 366138 508046 396678 508102
rect 396734 508046 396802 508102
rect 396858 508046 427398 508102
rect 427454 508046 427522 508102
rect 427578 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 474518 508102
rect 474574 508046 474642 508102
rect 474698 508046 505238 508102
rect 505294 508046 505362 508102
rect 505418 508046 535958 508102
rect 536014 508046 536082 508102
rect 536138 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 128394 507978
rect 128450 507922 128518 507978
rect 128574 507922 128642 507978
rect 128698 507922 128766 507978
rect 128822 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 164518 507978
rect 164574 507922 164642 507978
rect 164698 507922 195238 507978
rect 195294 507922 195362 507978
rect 195418 507922 220554 507978
rect 220610 507922 220678 507978
rect 220734 507922 220802 507978
rect 220858 507922 220926 507978
rect 220982 507922 251274 507978
rect 251330 507922 251398 507978
rect 251454 507922 251522 507978
rect 251578 507922 251646 507978
rect 251702 507922 281994 507978
rect 282050 507922 282118 507978
rect 282174 507922 282242 507978
rect 282298 507922 282366 507978
rect 282422 507922 304518 507978
rect 304574 507922 304642 507978
rect 304698 507922 335238 507978
rect 335294 507922 335362 507978
rect 335418 507922 365958 507978
rect 366014 507922 366082 507978
rect 366138 507922 396678 507978
rect 396734 507922 396802 507978
rect 396858 507922 427398 507978
rect 427454 507922 427522 507978
rect 427578 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 474518 507978
rect 474574 507922 474642 507978
rect 474698 507922 505238 507978
rect 505294 507922 505362 507978
rect 505418 507922 535958 507978
rect 536014 507922 536082 507978
rect 536138 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect 445996 499798 474980 499814
rect 445996 499742 446012 499798
rect 446068 499742 474908 499798
rect 474964 499742 474980 499798
rect 445996 499726 474980 499742
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496328 132114 496350
rect 40382 496294 67964 496328
rect -1916 496272 67964 496294
rect 68020 496272 68088 496328
rect 68144 496272 68212 496328
rect 68268 496272 68336 496328
rect 68392 496272 68460 496328
rect 68516 496272 68584 496328
rect 68640 496272 68708 496328
rect 68764 496272 68832 496328
rect 68888 496272 68956 496328
rect 69012 496272 69080 496328
rect 69136 496272 69204 496328
rect 69260 496272 69328 496328
rect 69384 496272 69452 496328
rect 69508 496272 69576 496328
rect 69632 496272 69700 496328
rect 69756 496272 69824 496328
rect 69880 496272 69948 496328
rect 70004 496272 70072 496328
rect 70128 496272 70196 496328
rect 70252 496272 70320 496328
rect 70376 496272 70444 496328
rect 70500 496272 70568 496328
rect 70624 496272 70692 496328
rect 70748 496272 70816 496328
rect 70872 496272 70940 496328
rect 70996 496272 71064 496328
rect 71120 496272 71188 496328
rect 71244 496272 71312 496328
rect 71368 496272 71436 496328
rect 71492 496272 71560 496328
rect 71616 496272 71684 496328
rect 71740 496272 71808 496328
rect 71864 496272 71932 496328
rect 71988 496272 72056 496328
rect 72112 496272 72180 496328
rect 72236 496272 72304 496328
rect 72360 496272 72428 496328
rect 72484 496272 72552 496328
rect 72608 496272 72676 496328
rect 72732 496272 72800 496328
rect 72856 496272 72924 496328
rect 72980 496272 73048 496328
rect 73104 496272 73172 496328
rect 73228 496272 73296 496328
rect 73352 496272 73420 496328
rect 73476 496272 73544 496328
rect 73600 496272 73668 496328
rect 73724 496272 73792 496328
rect 73848 496272 73916 496328
rect 73972 496272 74040 496328
rect 74096 496272 74164 496328
rect 74220 496272 74288 496328
rect 74344 496272 74412 496328
rect 74468 496272 74536 496328
rect 74592 496272 74660 496328
rect 74716 496294 132114 496328
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 224274 496350
rect 224330 496294 224398 496350
rect 224454 496294 224522 496350
rect 224578 496294 224646 496350
rect 224702 496294 254994 496350
rect 255050 496294 255118 496350
rect 255174 496294 255242 496350
rect 255298 496294 255366 496350
rect 255422 496294 285714 496350
rect 285770 496294 285838 496350
rect 285894 496294 285962 496350
rect 286018 496294 286086 496350
rect 286142 496294 319878 496350
rect 319934 496294 320002 496350
rect 320058 496294 350598 496350
rect 350654 496294 350722 496350
rect 350778 496294 381318 496350
rect 381374 496294 381442 496350
rect 381498 496294 412038 496350
rect 412094 496294 412162 496350
rect 412218 496294 442758 496350
rect 442814 496294 442882 496350
rect 442938 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 489878 496350
rect 489934 496294 490002 496350
rect 490058 496294 520598 496350
rect 520654 496294 520722 496350
rect 520778 496294 551318 496350
rect 551374 496294 551442 496350
rect 551498 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 74716 496272 597980 496294
rect -1916 496226 597980 496272
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 224274 496226
rect 224330 496170 224398 496226
rect 224454 496170 224522 496226
rect 224578 496170 224646 496226
rect 224702 496170 254994 496226
rect 255050 496170 255118 496226
rect 255174 496170 255242 496226
rect 255298 496170 255366 496226
rect 255422 496170 285714 496226
rect 285770 496170 285838 496226
rect 285894 496170 285962 496226
rect 286018 496170 286086 496226
rect 286142 496170 319878 496226
rect 319934 496170 320002 496226
rect 320058 496170 350598 496226
rect 350654 496170 350722 496226
rect 350778 496170 381318 496226
rect 381374 496170 381442 496226
rect 381498 496170 412038 496226
rect 412094 496170 412162 496226
rect 412218 496170 442758 496226
rect 442814 496170 442882 496226
rect 442938 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 489878 496226
rect 489934 496170 490002 496226
rect 490058 496170 520598 496226
rect 520654 496170 520722 496226
rect 520778 496170 551318 496226
rect 551374 496170 551442 496226
rect 551498 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496088 132114 496102
rect 40382 496046 68208 496088
rect -1916 496032 68208 496046
rect 68264 496032 68332 496088
rect 68388 496032 68456 496088
rect 68512 496032 68580 496088
rect 68636 496032 68704 496088
rect 68760 496032 68828 496088
rect 68884 496032 68952 496088
rect 69008 496032 69076 496088
rect 69132 496032 69200 496088
rect 69256 496032 69324 496088
rect 69380 496032 69448 496088
rect 69504 496032 69572 496088
rect 69628 496032 69696 496088
rect 69752 496032 69820 496088
rect 69876 496032 69944 496088
rect 70000 496032 70068 496088
rect 70124 496032 70192 496088
rect 70248 496032 70316 496088
rect 70372 496032 70440 496088
rect 70496 496032 70564 496088
rect 70620 496032 70688 496088
rect 70744 496032 70812 496088
rect 70868 496032 70936 496088
rect 70992 496032 71060 496088
rect 71116 496032 71184 496088
rect 71240 496032 71308 496088
rect 71364 496032 71432 496088
rect 71488 496032 71556 496088
rect 71612 496032 71680 496088
rect 71736 496032 71804 496088
rect 71860 496032 71928 496088
rect 71984 496032 72052 496088
rect 72108 496032 72176 496088
rect 72232 496032 72300 496088
rect 72356 496032 72424 496088
rect 72480 496032 72548 496088
rect 72604 496032 72672 496088
rect 72728 496032 72796 496088
rect 72852 496032 72920 496088
rect 72976 496032 73044 496088
rect 73100 496032 73168 496088
rect 73224 496032 73292 496088
rect 73348 496032 73416 496088
rect 73472 496032 73540 496088
rect 73596 496032 73664 496088
rect 73720 496032 73788 496088
rect 73844 496032 73912 496088
rect 73968 496032 74036 496088
rect 74092 496032 74160 496088
rect 74216 496032 74284 496088
rect 74340 496032 74408 496088
rect 74464 496032 74532 496088
rect 74588 496032 74656 496088
rect 74712 496046 132114 496088
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 224274 496102
rect 224330 496046 224398 496102
rect 224454 496046 224522 496102
rect 224578 496046 224646 496102
rect 224702 496046 254994 496102
rect 255050 496046 255118 496102
rect 255174 496046 255242 496102
rect 255298 496046 255366 496102
rect 255422 496046 285714 496102
rect 285770 496046 285838 496102
rect 285894 496046 285962 496102
rect 286018 496046 286086 496102
rect 286142 496046 319878 496102
rect 319934 496046 320002 496102
rect 320058 496046 350598 496102
rect 350654 496046 350722 496102
rect 350778 496046 381318 496102
rect 381374 496046 381442 496102
rect 381498 496046 412038 496102
rect 412094 496046 412162 496102
rect 412218 496046 442758 496102
rect 442814 496046 442882 496102
rect 442938 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 489878 496102
rect 489934 496046 490002 496102
rect 490058 496046 520598 496102
rect 520654 496046 520722 496102
rect 520778 496046 551318 496102
rect 551374 496046 551442 496102
rect 551498 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 74712 496032 597980 496046
rect -1916 495978 597980 496032
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 132114 495978
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 224274 495978
rect 224330 495922 224398 495978
rect 224454 495922 224522 495978
rect 224578 495922 224646 495978
rect 224702 495922 254994 495978
rect 255050 495922 255118 495978
rect 255174 495922 255242 495978
rect 255298 495922 255366 495978
rect 255422 495922 285714 495978
rect 285770 495922 285838 495978
rect 285894 495922 285962 495978
rect 286018 495922 286086 495978
rect 286142 495922 319878 495978
rect 319934 495922 320002 495978
rect 320058 495922 350598 495978
rect 350654 495922 350722 495978
rect 350778 495922 381318 495978
rect 381374 495922 381442 495978
rect 381498 495922 412038 495978
rect 412094 495922 412162 495978
rect 412218 495922 442758 495978
rect 442814 495922 442882 495978
rect 442938 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 489878 495978
rect 489934 495922 490002 495978
rect 490058 495922 520598 495978
rect 520654 495922 520722 495978
rect 520778 495922 551318 495978
rect 551374 495922 551442 495978
rect 551498 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 66954 490350
rect 67010 490294 67078 490350
rect 67134 490294 67202 490350
rect 67258 490294 67326 490350
rect 67382 490294 97674 490350
rect 97730 490294 97798 490350
rect 97854 490294 97922 490350
rect 97978 490294 98046 490350
rect 98102 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 220554 490350
rect 220610 490294 220678 490350
rect 220734 490294 220802 490350
rect 220858 490294 220926 490350
rect 220982 490294 251274 490350
rect 251330 490294 251398 490350
rect 251454 490294 251522 490350
rect 251578 490294 251646 490350
rect 251702 490294 281994 490350
rect 282050 490294 282118 490350
rect 282174 490294 282242 490350
rect 282298 490294 282366 490350
rect 282422 490294 304518 490350
rect 304574 490294 304642 490350
rect 304698 490294 335238 490350
rect 335294 490294 335362 490350
rect 335418 490294 365958 490350
rect 366014 490294 366082 490350
rect 366138 490294 396678 490350
rect 396734 490294 396802 490350
rect 396858 490294 427398 490350
rect 427454 490294 427522 490350
rect 427578 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 474518 490350
rect 474574 490294 474642 490350
rect 474698 490294 505238 490350
rect 505294 490294 505362 490350
rect 505418 490294 535958 490350
rect 536014 490294 536082 490350
rect 536138 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 66954 490226
rect 67010 490170 67078 490226
rect 67134 490170 67202 490226
rect 67258 490170 67326 490226
rect 67382 490170 97674 490226
rect 97730 490170 97798 490226
rect 97854 490170 97922 490226
rect 97978 490170 98046 490226
rect 98102 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 220554 490226
rect 220610 490170 220678 490226
rect 220734 490170 220802 490226
rect 220858 490170 220926 490226
rect 220982 490170 251274 490226
rect 251330 490170 251398 490226
rect 251454 490170 251522 490226
rect 251578 490170 251646 490226
rect 251702 490170 281994 490226
rect 282050 490170 282118 490226
rect 282174 490170 282242 490226
rect 282298 490170 282366 490226
rect 282422 490170 304518 490226
rect 304574 490170 304642 490226
rect 304698 490170 335238 490226
rect 335294 490170 335362 490226
rect 335418 490170 365958 490226
rect 366014 490170 366082 490226
rect 366138 490170 396678 490226
rect 396734 490170 396802 490226
rect 396858 490170 427398 490226
rect 427454 490170 427522 490226
rect 427578 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 474518 490226
rect 474574 490170 474642 490226
rect 474698 490170 505238 490226
rect 505294 490170 505362 490226
rect 505418 490170 535958 490226
rect 536014 490170 536082 490226
rect 536138 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 66954 490102
rect 67010 490046 67078 490102
rect 67134 490046 67202 490102
rect 67258 490046 67326 490102
rect 67382 490046 97674 490102
rect 97730 490046 97798 490102
rect 97854 490046 97922 490102
rect 97978 490046 98046 490102
rect 98102 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 220554 490102
rect 220610 490046 220678 490102
rect 220734 490046 220802 490102
rect 220858 490046 220926 490102
rect 220982 490046 251274 490102
rect 251330 490046 251398 490102
rect 251454 490046 251522 490102
rect 251578 490046 251646 490102
rect 251702 490046 281994 490102
rect 282050 490046 282118 490102
rect 282174 490046 282242 490102
rect 282298 490046 282366 490102
rect 282422 490046 304518 490102
rect 304574 490046 304642 490102
rect 304698 490046 335238 490102
rect 335294 490046 335362 490102
rect 335418 490046 365958 490102
rect 366014 490046 366082 490102
rect 366138 490046 396678 490102
rect 396734 490046 396802 490102
rect 396858 490046 427398 490102
rect 427454 490046 427522 490102
rect 427578 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 474518 490102
rect 474574 490046 474642 490102
rect 474698 490046 505238 490102
rect 505294 490046 505362 490102
rect 505418 490046 535958 490102
rect 536014 490046 536082 490102
rect 536138 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 66954 489978
rect 67010 489922 67078 489978
rect 67134 489922 67202 489978
rect 67258 489922 67326 489978
rect 67382 489922 97674 489978
rect 97730 489922 97798 489978
rect 97854 489922 97922 489978
rect 97978 489922 98046 489978
rect 98102 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 220554 489978
rect 220610 489922 220678 489978
rect 220734 489922 220802 489978
rect 220858 489922 220926 489978
rect 220982 489922 251274 489978
rect 251330 489922 251398 489978
rect 251454 489922 251522 489978
rect 251578 489922 251646 489978
rect 251702 489922 281994 489978
rect 282050 489922 282118 489978
rect 282174 489922 282242 489978
rect 282298 489922 282366 489978
rect 282422 489922 304518 489978
rect 304574 489922 304642 489978
rect 304698 489922 335238 489978
rect 335294 489922 335362 489978
rect 335418 489922 365958 489978
rect 366014 489922 366082 489978
rect 366138 489922 396678 489978
rect 396734 489922 396802 489978
rect 396858 489922 427398 489978
rect 427454 489922 427522 489978
rect 427578 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 474518 489978
rect 474574 489922 474642 489978
rect 474698 489922 505238 489978
rect 505294 489922 505362 489978
rect 505418 489922 535958 489978
rect 536014 489922 536082 489978
rect 536138 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect 169580 488098 303396 488114
rect 169580 488042 169596 488098
rect 169652 488042 303324 488098
rect 303380 488042 303396 488098
rect 169580 488026 303396 488042
rect 166220 479638 303508 479654
rect 166220 479582 166236 479638
rect 166292 479582 303436 479638
rect 303492 479582 303508 479638
rect 166220 479566 303508 479582
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 101394 478350
rect 101450 478294 101518 478350
rect 101574 478294 101642 478350
rect 101698 478294 101766 478350
rect 101822 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 224274 478350
rect 224330 478294 224398 478350
rect 224454 478294 224522 478350
rect 224578 478294 224646 478350
rect 224702 478294 254994 478350
rect 255050 478294 255118 478350
rect 255174 478294 255242 478350
rect 255298 478294 255366 478350
rect 255422 478294 285714 478350
rect 285770 478294 285838 478350
rect 285894 478294 285962 478350
rect 286018 478294 286086 478350
rect 286142 478294 319878 478350
rect 319934 478294 320002 478350
rect 320058 478294 350598 478350
rect 350654 478294 350722 478350
rect 350778 478294 381318 478350
rect 381374 478294 381442 478350
rect 381498 478294 412038 478350
rect 412094 478294 412162 478350
rect 412218 478294 442758 478350
rect 442814 478294 442882 478350
rect 442938 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 489878 478350
rect 489934 478294 490002 478350
rect 490058 478294 520598 478350
rect 520654 478294 520722 478350
rect 520778 478294 551318 478350
rect 551374 478294 551442 478350
rect 551498 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 101394 478226
rect 101450 478170 101518 478226
rect 101574 478170 101642 478226
rect 101698 478170 101766 478226
rect 101822 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 224274 478226
rect 224330 478170 224398 478226
rect 224454 478170 224522 478226
rect 224578 478170 224646 478226
rect 224702 478170 254994 478226
rect 255050 478170 255118 478226
rect 255174 478170 255242 478226
rect 255298 478170 255366 478226
rect 255422 478170 285714 478226
rect 285770 478170 285838 478226
rect 285894 478170 285962 478226
rect 286018 478170 286086 478226
rect 286142 478170 319878 478226
rect 319934 478170 320002 478226
rect 320058 478170 350598 478226
rect 350654 478170 350722 478226
rect 350778 478170 381318 478226
rect 381374 478170 381442 478226
rect 381498 478170 412038 478226
rect 412094 478170 412162 478226
rect 412218 478170 442758 478226
rect 442814 478170 442882 478226
rect 442938 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 489878 478226
rect 489934 478170 490002 478226
rect 490058 478170 520598 478226
rect 520654 478170 520722 478226
rect 520778 478170 551318 478226
rect 551374 478170 551442 478226
rect 551498 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 101394 478102
rect 101450 478046 101518 478102
rect 101574 478046 101642 478102
rect 101698 478046 101766 478102
rect 101822 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 224274 478102
rect 224330 478046 224398 478102
rect 224454 478046 224522 478102
rect 224578 478046 224646 478102
rect 224702 478046 254994 478102
rect 255050 478046 255118 478102
rect 255174 478046 255242 478102
rect 255298 478046 255366 478102
rect 255422 478046 285714 478102
rect 285770 478046 285838 478102
rect 285894 478046 285962 478102
rect 286018 478046 286086 478102
rect 286142 478046 319878 478102
rect 319934 478046 320002 478102
rect 320058 478046 350598 478102
rect 350654 478046 350722 478102
rect 350778 478046 381318 478102
rect 381374 478046 381442 478102
rect 381498 478046 412038 478102
rect 412094 478046 412162 478102
rect 412218 478046 442758 478102
rect 442814 478046 442882 478102
rect 442938 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 489878 478102
rect 489934 478046 490002 478102
rect 490058 478046 520598 478102
rect 520654 478046 520722 478102
rect 520778 478046 551318 478102
rect 551374 478046 551442 478102
rect 551498 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 101394 477978
rect 101450 477922 101518 477978
rect 101574 477922 101642 477978
rect 101698 477922 101766 477978
rect 101822 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 224274 477978
rect 224330 477922 224398 477978
rect 224454 477922 224522 477978
rect 224578 477922 224646 477978
rect 224702 477922 254994 477978
rect 255050 477922 255118 477978
rect 255174 477922 255242 477978
rect 255298 477922 255366 477978
rect 255422 477922 285714 477978
rect 285770 477922 285838 477978
rect 285894 477922 285962 477978
rect 286018 477922 286086 477978
rect 286142 477922 319878 477978
rect 319934 477922 320002 477978
rect 320058 477922 350598 477978
rect 350654 477922 350722 477978
rect 350778 477922 381318 477978
rect 381374 477922 381442 477978
rect 381498 477922 412038 477978
rect 412094 477922 412162 477978
rect 412218 477922 442758 477978
rect 442814 477922 442882 477978
rect 442938 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 489878 477978
rect 489934 477922 490002 477978
rect 490058 477922 520598 477978
rect 520654 477922 520722 477978
rect 520778 477922 551318 477978
rect 551374 477922 551442 477978
rect 551498 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect 164540 472618 303284 472634
rect 164540 472562 164556 472618
rect 164612 472562 303212 472618
rect 303268 472562 303284 472618
rect 164540 472546 303284 472562
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 220554 472350
rect 220610 472294 220678 472350
rect 220734 472294 220802 472350
rect 220858 472294 220926 472350
rect 220982 472294 251274 472350
rect 251330 472294 251398 472350
rect 251454 472294 251522 472350
rect 251578 472294 251646 472350
rect 251702 472294 281994 472350
rect 282050 472294 282118 472350
rect 282174 472294 282242 472350
rect 282298 472294 282366 472350
rect 282422 472294 304518 472350
rect 304574 472294 304642 472350
rect 304698 472294 335238 472350
rect 335294 472294 335362 472350
rect 335418 472294 365958 472350
rect 366014 472294 366082 472350
rect 366138 472294 396678 472350
rect 396734 472294 396802 472350
rect 396858 472294 427398 472350
rect 427454 472294 427522 472350
rect 427578 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 474518 472350
rect 474574 472294 474642 472350
rect 474698 472294 505238 472350
rect 505294 472294 505362 472350
rect 505418 472294 535958 472350
rect 536014 472294 536082 472350
rect 536138 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 220554 472226
rect 220610 472170 220678 472226
rect 220734 472170 220802 472226
rect 220858 472170 220926 472226
rect 220982 472170 251274 472226
rect 251330 472170 251398 472226
rect 251454 472170 251522 472226
rect 251578 472170 251646 472226
rect 251702 472170 281994 472226
rect 282050 472170 282118 472226
rect 282174 472170 282242 472226
rect 282298 472170 282366 472226
rect 282422 472170 304518 472226
rect 304574 472170 304642 472226
rect 304698 472170 335238 472226
rect 335294 472170 335362 472226
rect 335418 472170 365958 472226
rect 366014 472170 366082 472226
rect 366138 472170 396678 472226
rect 396734 472170 396802 472226
rect 396858 472170 427398 472226
rect 427454 472170 427522 472226
rect 427578 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 474518 472226
rect 474574 472170 474642 472226
rect 474698 472170 505238 472226
rect 505294 472170 505362 472226
rect 505418 472170 535958 472226
rect 536014 472170 536082 472226
rect 536138 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 220554 472102
rect 220610 472046 220678 472102
rect 220734 472046 220802 472102
rect 220858 472046 220926 472102
rect 220982 472046 251274 472102
rect 251330 472046 251398 472102
rect 251454 472046 251522 472102
rect 251578 472046 251646 472102
rect 251702 472046 281994 472102
rect 282050 472046 282118 472102
rect 282174 472046 282242 472102
rect 282298 472046 282366 472102
rect 282422 472046 304518 472102
rect 304574 472046 304642 472102
rect 304698 472046 335238 472102
rect 335294 472046 335362 472102
rect 335418 472046 365958 472102
rect 366014 472046 366082 472102
rect 366138 472046 396678 472102
rect 396734 472046 396802 472102
rect 396858 472046 427398 472102
rect 427454 472046 427522 472102
rect 427578 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 474518 472102
rect 474574 472046 474642 472102
rect 474698 472046 505238 472102
rect 505294 472046 505362 472102
rect 505418 472046 535958 472102
rect 536014 472046 536082 472102
rect 536138 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 220554 471978
rect 220610 471922 220678 471978
rect 220734 471922 220802 471978
rect 220858 471922 220926 471978
rect 220982 471922 251274 471978
rect 251330 471922 251398 471978
rect 251454 471922 251522 471978
rect 251578 471922 251646 471978
rect 251702 471922 281994 471978
rect 282050 471922 282118 471978
rect 282174 471922 282242 471978
rect 282298 471922 282366 471978
rect 282422 471922 304518 471978
rect 304574 471922 304642 471978
rect 304698 471922 335238 471978
rect 335294 471922 335362 471978
rect 335418 471922 365958 471978
rect 366014 471922 366082 471978
rect 366138 471922 396678 471978
rect 396734 471922 396802 471978
rect 396858 471922 427398 471978
rect 427454 471922 427522 471978
rect 427578 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 474518 471978
rect 474574 471922 474642 471978
rect 474698 471922 505238 471978
rect 505294 471922 505362 471978
rect 505418 471922 535958 471978
rect 536014 471922 536082 471978
rect 536138 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 224274 460350
rect 224330 460294 224398 460350
rect 224454 460294 224522 460350
rect 224578 460294 224646 460350
rect 224702 460294 254994 460350
rect 255050 460294 255118 460350
rect 255174 460294 255242 460350
rect 255298 460294 255366 460350
rect 255422 460294 285714 460350
rect 285770 460294 285838 460350
rect 285894 460294 285962 460350
rect 286018 460294 286086 460350
rect 286142 460294 319878 460350
rect 319934 460294 320002 460350
rect 320058 460294 350598 460350
rect 350654 460294 350722 460350
rect 350778 460294 381318 460350
rect 381374 460294 381442 460350
rect 381498 460294 412038 460350
rect 412094 460294 412162 460350
rect 412218 460294 442758 460350
rect 442814 460294 442882 460350
rect 442938 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 489878 460350
rect 489934 460294 490002 460350
rect 490058 460294 520598 460350
rect 520654 460294 520722 460350
rect 520778 460294 551318 460350
rect 551374 460294 551442 460350
rect 551498 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 224274 460226
rect 224330 460170 224398 460226
rect 224454 460170 224522 460226
rect 224578 460170 224646 460226
rect 224702 460170 254994 460226
rect 255050 460170 255118 460226
rect 255174 460170 255242 460226
rect 255298 460170 255366 460226
rect 255422 460170 285714 460226
rect 285770 460170 285838 460226
rect 285894 460170 285962 460226
rect 286018 460170 286086 460226
rect 286142 460170 319878 460226
rect 319934 460170 320002 460226
rect 320058 460170 350598 460226
rect 350654 460170 350722 460226
rect 350778 460170 381318 460226
rect 381374 460170 381442 460226
rect 381498 460170 412038 460226
rect 412094 460170 412162 460226
rect 412218 460170 442758 460226
rect 442814 460170 442882 460226
rect 442938 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 489878 460226
rect 489934 460170 490002 460226
rect 490058 460170 520598 460226
rect 520654 460170 520722 460226
rect 520778 460170 551318 460226
rect 551374 460170 551442 460226
rect 551498 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 224274 460102
rect 224330 460046 224398 460102
rect 224454 460046 224522 460102
rect 224578 460046 224646 460102
rect 224702 460046 254994 460102
rect 255050 460046 255118 460102
rect 255174 460046 255242 460102
rect 255298 460046 255366 460102
rect 255422 460046 285714 460102
rect 285770 460046 285838 460102
rect 285894 460046 285962 460102
rect 286018 460046 286086 460102
rect 286142 460046 319878 460102
rect 319934 460046 320002 460102
rect 320058 460046 350598 460102
rect 350654 460046 350722 460102
rect 350778 460046 381318 460102
rect 381374 460046 381442 460102
rect 381498 460046 412038 460102
rect 412094 460046 412162 460102
rect 412218 460046 442758 460102
rect 442814 460046 442882 460102
rect 442938 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 489878 460102
rect 489934 460046 490002 460102
rect 490058 460046 520598 460102
rect 520654 460046 520722 460102
rect 520778 460046 551318 460102
rect 551374 460046 551442 460102
rect 551498 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 224274 459978
rect 224330 459922 224398 459978
rect 224454 459922 224522 459978
rect 224578 459922 224646 459978
rect 224702 459922 254994 459978
rect 255050 459922 255118 459978
rect 255174 459922 255242 459978
rect 255298 459922 255366 459978
rect 255422 459922 285714 459978
rect 285770 459922 285838 459978
rect 285894 459922 285962 459978
rect 286018 459922 286086 459978
rect 286142 459922 319878 459978
rect 319934 459922 320002 459978
rect 320058 459922 350598 459978
rect 350654 459922 350722 459978
rect 350778 459922 381318 459978
rect 381374 459922 381442 459978
rect 381498 459922 412038 459978
rect 412094 459922 412162 459978
rect 412218 459922 442758 459978
rect 442814 459922 442882 459978
rect 442938 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 489878 459978
rect 489934 459922 490002 459978
rect 490058 459922 520598 459978
rect 520654 459922 520722 459978
rect 520778 459922 551318 459978
rect 551374 459922 551442 459978
rect 551498 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 220554 454350
rect 220610 454294 220678 454350
rect 220734 454294 220802 454350
rect 220858 454294 220926 454350
rect 220982 454294 251274 454350
rect 251330 454294 251398 454350
rect 251454 454294 251522 454350
rect 251578 454294 251646 454350
rect 251702 454294 281994 454350
rect 282050 454294 282118 454350
rect 282174 454294 282242 454350
rect 282298 454294 282366 454350
rect 282422 454294 304518 454350
rect 304574 454294 304642 454350
rect 304698 454294 335238 454350
rect 335294 454294 335362 454350
rect 335418 454294 365958 454350
rect 366014 454294 366082 454350
rect 366138 454294 396678 454350
rect 396734 454294 396802 454350
rect 396858 454294 427398 454350
rect 427454 454294 427522 454350
rect 427578 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 474518 454350
rect 474574 454294 474642 454350
rect 474698 454294 505238 454350
rect 505294 454294 505362 454350
rect 505418 454294 535958 454350
rect 536014 454294 536082 454350
rect 536138 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 220554 454226
rect 220610 454170 220678 454226
rect 220734 454170 220802 454226
rect 220858 454170 220926 454226
rect 220982 454170 251274 454226
rect 251330 454170 251398 454226
rect 251454 454170 251522 454226
rect 251578 454170 251646 454226
rect 251702 454170 281994 454226
rect 282050 454170 282118 454226
rect 282174 454170 282242 454226
rect 282298 454170 282366 454226
rect 282422 454170 304518 454226
rect 304574 454170 304642 454226
rect 304698 454170 335238 454226
rect 335294 454170 335362 454226
rect 335418 454170 365958 454226
rect 366014 454170 366082 454226
rect 366138 454170 396678 454226
rect 396734 454170 396802 454226
rect 396858 454170 427398 454226
rect 427454 454170 427522 454226
rect 427578 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 474518 454226
rect 474574 454170 474642 454226
rect 474698 454170 505238 454226
rect 505294 454170 505362 454226
rect 505418 454170 535958 454226
rect 536014 454170 536082 454226
rect 536138 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 220554 454102
rect 220610 454046 220678 454102
rect 220734 454046 220802 454102
rect 220858 454046 220926 454102
rect 220982 454046 251274 454102
rect 251330 454046 251398 454102
rect 251454 454046 251522 454102
rect 251578 454046 251646 454102
rect 251702 454046 281994 454102
rect 282050 454046 282118 454102
rect 282174 454046 282242 454102
rect 282298 454046 282366 454102
rect 282422 454046 304518 454102
rect 304574 454046 304642 454102
rect 304698 454046 335238 454102
rect 335294 454046 335362 454102
rect 335418 454046 365958 454102
rect 366014 454046 366082 454102
rect 366138 454046 396678 454102
rect 396734 454046 396802 454102
rect 396858 454046 427398 454102
rect 427454 454046 427522 454102
rect 427578 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 474518 454102
rect 474574 454046 474642 454102
rect 474698 454046 505238 454102
rect 505294 454046 505362 454102
rect 505418 454046 535958 454102
rect 536014 454046 536082 454102
rect 536138 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 220554 453978
rect 220610 453922 220678 453978
rect 220734 453922 220802 453978
rect 220858 453922 220926 453978
rect 220982 453922 251274 453978
rect 251330 453922 251398 453978
rect 251454 453922 251522 453978
rect 251578 453922 251646 453978
rect 251702 453922 281994 453978
rect 282050 453922 282118 453978
rect 282174 453922 282242 453978
rect 282298 453922 282366 453978
rect 282422 453922 304518 453978
rect 304574 453922 304642 453978
rect 304698 453922 335238 453978
rect 335294 453922 335362 453978
rect 335418 453922 365958 453978
rect 366014 453922 366082 453978
rect 366138 453922 396678 453978
rect 396734 453922 396802 453978
rect 396858 453922 427398 453978
rect 427454 453922 427522 453978
rect 427578 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 474518 453978
rect 474574 453922 474642 453978
rect 474698 453922 505238 453978
rect 505294 453922 505362 453978
rect 505418 453922 535958 453978
rect 536014 453922 536082 453978
rect 536138 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect 478028 451018 590788 451034
rect 478028 450962 478044 451018
rect 478100 450962 590716 451018
rect 590772 450962 590788 451018
rect 478028 450946 590788 450962
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 224274 442350
rect 224330 442294 224398 442350
rect 224454 442294 224522 442350
rect 224578 442294 224646 442350
rect 224702 442294 254994 442350
rect 255050 442294 255118 442350
rect 255174 442294 255242 442350
rect 255298 442294 255366 442350
rect 255422 442294 285714 442350
rect 285770 442294 285838 442350
rect 285894 442294 285962 442350
rect 286018 442294 286086 442350
rect 286142 442294 319878 442350
rect 319934 442294 320002 442350
rect 320058 442294 350598 442350
rect 350654 442294 350722 442350
rect 350778 442294 381318 442350
rect 381374 442294 381442 442350
rect 381498 442294 412038 442350
rect 412094 442294 412162 442350
rect 412218 442294 442758 442350
rect 442814 442294 442882 442350
rect 442938 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 224274 442226
rect 224330 442170 224398 442226
rect 224454 442170 224522 442226
rect 224578 442170 224646 442226
rect 224702 442170 254994 442226
rect 255050 442170 255118 442226
rect 255174 442170 255242 442226
rect 255298 442170 255366 442226
rect 255422 442170 285714 442226
rect 285770 442170 285838 442226
rect 285894 442170 285962 442226
rect 286018 442170 286086 442226
rect 286142 442170 319878 442226
rect 319934 442170 320002 442226
rect 320058 442170 350598 442226
rect 350654 442170 350722 442226
rect 350778 442170 381318 442226
rect 381374 442170 381442 442226
rect 381498 442170 412038 442226
rect 412094 442170 412162 442226
rect 412218 442170 442758 442226
rect 442814 442170 442882 442226
rect 442938 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 224274 442102
rect 224330 442046 224398 442102
rect 224454 442046 224522 442102
rect 224578 442046 224646 442102
rect 224702 442046 254994 442102
rect 255050 442046 255118 442102
rect 255174 442046 255242 442102
rect 255298 442046 255366 442102
rect 255422 442046 285714 442102
rect 285770 442046 285838 442102
rect 285894 442046 285962 442102
rect 286018 442046 286086 442102
rect 286142 442046 319878 442102
rect 319934 442046 320002 442102
rect 320058 442046 350598 442102
rect 350654 442046 350722 442102
rect 350778 442046 381318 442102
rect 381374 442046 381442 442102
rect 381498 442046 412038 442102
rect 412094 442046 412162 442102
rect 412218 442046 442758 442102
rect 442814 442046 442882 442102
rect 442938 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 224274 441978
rect 224330 441922 224398 441978
rect 224454 441922 224522 441978
rect 224578 441922 224646 441978
rect 224702 441922 254994 441978
rect 255050 441922 255118 441978
rect 255174 441922 255242 441978
rect 255298 441922 255366 441978
rect 255422 441922 285714 441978
rect 285770 441922 285838 441978
rect 285894 441922 285962 441978
rect 286018 441922 286086 441978
rect 286142 441922 319878 441978
rect 319934 441922 320002 441978
rect 320058 441922 350598 441978
rect 350654 441922 350722 441978
rect 350778 441922 381318 441978
rect 381374 441922 381442 441978
rect 381498 441922 412038 441978
rect 412094 441922 412162 441978
rect 412218 441922 442758 441978
rect 442814 441922 442882 441978
rect 442938 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 220554 436350
rect 220610 436294 220678 436350
rect 220734 436294 220802 436350
rect 220858 436294 220926 436350
rect 220982 436294 251274 436350
rect 251330 436294 251398 436350
rect 251454 436294 251522 436350
rect 251578 436294 251646 436350
rect 251702 436294 281994 436350
rect 282050 436294 282118 436350
rect 282174 436294 282242 436350
rect 282298 436294 282366 436350
rect 282422 436294 304518 436350
rect 304574 436294 304642 436350
rect 304698 436294 335238 436350
rect 335294 436294 335362 436350
rect 335418 436294 365958 436350
rect 366014 436294 366082 436350
rect 366138 436294 396678 436350
rect 396734 436294 396802 436350
rect 396858 436294 427398 436350
rect 427454 436294 427522 436350
rect 427578 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 220554 436226
rect 220610 436170 220678 436226
rect 220734 436170 220802 436226
rect 220858 436170 220926 436226
rect 220982 436170 251274 436226
rect 251330 436170 251398 436226
rect 251454 436170 251522 436226
rect 251578 436170 251646 436226
rect 251702 436170 281994 436226
rect 282050 436170 282118 436226
rect 282174 436170 282242 436226
rect 282298 436170 282366 436226
rect 282422 436170 304518 436226
rect 304574 436170 304642 436226
rect 304698 436170 335238 436226
rect 335294 436170 335362 436226
rect 335418 436170 365958 436226
rect 366014 436170 366082 436226
rect 366138 436170 396678 436226
rect 396734 436170 396802 436226
rect 396858 436170 427398 436226
rect 427454 436170 427522 436226
rect 427578 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 220554 436102
rect 220610 436046 220678 436102
rect 220734 436046 220802 436102
rect 220858 436046 220926 436102
rect 220982 436046 251274 436102
rect 251330 436046 251398 436102
rect 251454 436046 251522 436102
rect 251578 436046 251646 436102
rect 251702 436046 281994 436102
rect 282050 436046 282118 436102
rect 282174 436046 282242 436102
rect 282298 436046 282366 436102
rect 282422 436046 304518 436102
rect 304574 436046 304642 436102
rect 304698 436046 335238 436102
rect 335294 436046 335362 436102
rect 335418 436046 365958 436102
rect 366014 436046 366082 436102
rect 366138 436046 396678 436102
rect 396734 436046 396802 436102
rect 396858 436046 427398 436102
rect 427454 436046 427522 436102
rect 427578 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 220554 435978
rect 220610 435922 220678 435978
rect 220734 435922 220802 435978
rect 220858 435922 220926 435978
rect 220982 435922 251274 435978
rect 251330 435922 251398 435978
rect 251454 435922 251522 435978
rect 251578 435922 251646 435978
rect 251702 435922 281994 435978
rect 282050 435922 282118 435978
rect 282174 435922 282242 435978
rect 282298 435922 282366 435978
rect 282422 435922 304518 435978
rect 304574 435922 304642 435978
rect 304698 435922 335238 435978
rect 335294 435922 335362 435978
rect 335418 435922 365958 435978
rect 366014 435922 366082 435978
rect 366138 435922 396678 435978
rect 396734 435922 396802 435978
rect 396858 435922 427398 435978
rect 427454 435922 427522 435978
rect 427578 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect 452716 433378 512388 433394
rect 452716 433322 452732 433378
rect 452788 433322 512316 433378
rect 512372 433322 512388 433378
rect 452716 433306 512388 433322
rect 479820 432478 498948 432494
rect 479820 432422 479836 432478
rect 479892 432422 498876 432478
rect 498932 432422 498948 432478
rect 479820 432406 498948 432422
rect 479596 432298 502980 432314
rect 479596 432242 479612 432298
rect 479668 432242 502908 432298
rect 502964 432242 502980 432298
rect 479596 432226 502980 432242
rect 82892 432118 276404 432134
rect 82892 432062 82908 432118
rect 82964 432062 276332 432118
rect 276388 432062 276404 432118
rect 82892 432046 276404 432062
rect 480044 432118 519108 432134
rect 480044 432062 480060 432118
rect 480116 432062 519036 432118
rect 519092 432062 519108 432118
rect 480044 432046 519108 432062
rect 77516 431938 288276 431954
rect 77516 431882 77532 431938
rect 77588 431882 288204 431938
rect 288260 431882 288276 431938
rect 77516 431866 288276 431882
rect 477916 431938 523140 431954
rect 477916 431882 477932 431938
rect 477988 431882 523068 431938
rect 523124 431882 523140 431938
rect 477916 431866 523140 431882
rect 69452 431038 300036 431054
rect 69452 430982 69468 431038
rect 69524 430982 299964 431038
rect 300020 430982 300036 431038
rect 69452 430966 300036 430982
rect 4940 430858 296676 430874
rect 4940 430802 4956 430858
rect 5012 430802 296604 430858
rect 296660 430802 296676 430858
rect 4940 430786 296676 430802
rect 4156 430138 298244 430154
rect 4156 430082 4172 430138
rect 4228 430082 298172 430138
rect 298228 430082 298244 430138
rect 4156 430066 298244 430082
rect 74828 429418 284916 429434
rect 74828 429362 74844 429418
rect 74900 429362 284844 429418
rect 284900 429362 284916 429418
rect 74828 429346 284916 429362
rect 80204 428518 298580 428534
rect 80204 428462 80220 428518
rect 80276 428462 298508 428518
rect 298564 428462 298580 428518
rect 80204 428446 298580 428462
rect 300844 427438 301604 427454
rect 300844 427382 300860 427438
rect 300916 427382 301532 427438
rect 301588 427382 301604 427438
rect 300844 427366 301604 427382
rect 56572 427258 281444 427274
rect 56572 427202 56588 427258
rect 56644 427202 281372 427258
rect 281428 427202 281444 427258
rect 56572 427186 281444 427202
rect 57020 427078 289844 427094
rect 57020 427022 57036 427078
rect 57092 427022 289772 427078
rect 289828 427022 289844 427078
rect 57020 427006 289844 427022
rect 4268 426898 298132 426914
rect 4268 426842 4284 426898
rect 4340 426842 298060 426898
rect 298116 426842 298132 426898
rect 4268 426826 298132 426842
rect 83116 425458 294884 425474
rect 83116 425402 83132 425458
rect 83188 425402 294812 425458
rect 294868 425402 294884 425458
rect 83116 425386 294884 425402
rect 83452 425278 301044 425294
rect 83452 425222 83468 425278
rect 83524 425222 300972 425278
rect 301028 425222 301044 425278
rect 83452 425206 301044 425222
rect 56684 425098 299924 425114
rect 56684 425042 56700 425098
rect 56756 425042 299852 425098
rect 299908 425042 299924 425098
rect 56684 425026 299924 425042
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 79878 424350
rect 79934 424294 80002 424350
rect 80058 424294 110598 424350
rect 110654 424294 110722 424350
rect 110778 424294 141318 424350
rect 141374 424294 141442 424350
rect 141498 424294 172038 424350
rect 172094 424294 172162 424350
rect 172218 424294 202758 424350
rect 202814 424294 202882 424350
rect 202938 424294 233478 424350
rect 233534 424294 233602 424350
rect 233658 424294 264198 424350
rect 264254 424294 264322 424350
rect 264378 424294 285714 424350
rect 285770 424294 285838 424350
rect 285894 424294 285962 424350
rect 286018 424294 286086 424350
rect 286142 424294 319878 424350
rect 319934 424294 320002 424350
rect 320058 424294 350598 424350
rect 350654 424294 350722 424350
rect 350778 424294 381318 424350
rect 381374 424294 381442 424350
rect 381498 424294 412038 424350
rect 412094 424294 412162 424350
rect 412218 424294 442758 424350
rect 442814 424294 442882 424350
rect 442938 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 499878 424350
rect 499934 424294 500002 424350
rect 500058 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 79878 424226
rect 79934 424170 80002 424226
rect 80058 424170 110598 424226
rect 110654 424170 110722 424226
rect 110778 424170 141318 424226
rect 141374 424170 141442 424226
rect 141498 424170 172038 424226
rect 172094 424170 172162 424226
rect 172218 424170 202758 424226
rect 202814 424170 202882 424226
rect 202938 424170 233478 424226
rect 233534 424170 233602 424226
rect 233658 424170 264198 424226
rect 264254 424170 264322 424226
rect 264378 424170 285714 424226
rect 285770 424170 285838 424226
rect 285894 424170 285962 424226
rect 286018 424170 286086 424226
rect 286142 424170 319878 424226
rect 319934 424170 320002 424226
rect 320058 424170 350598 424226
rect 350654 424170 350722 424226
rect 350778 424170 381318 424226
rect 381374 424170 381442 424226
rect 381498 424170 412038 424226
rect 412094 424170 412162 424226
rect 412218 424170 442758 424226
rect 442814 424170 442882 424226
rect 442938 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 499878 424226
rect 499934 424170 500002 424226
rect 500058 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 79878 424102
rect 79934 424046 80002 424102
rect 80058 424046 110598 424102
rect 110654 424046 110722 424102
rect 110778 424046 141318 424102
rect 141374 424046 141442 424102
rect 141498 424046 172038 424102
rect 172094 424046 172162 424102
rect 172218 424046 202758 424102
rect 202814 424046 202882 424102
rect 202938 424046 233478 424102
rect 233534 424046 233602 424102
rect 233658 424046 264198 424102
rect 264254 424046 264322 424102
rect 264378 424046 285714 424102
rect 285770 424046 285838 424102
rect 285894 424046 285962 424102
rect 286018 424046 286086 424102
rect 286142 424046 319878 424102
rect 319934 424046 320002 424102
rect 320058 424046 350598 424102
rect 350654 424046 350722 424102
rect 350778 424046 381318 424102
rect 381374 424046 381442 424102
rect 381498 424046 412038 424102
rect 412094 424046 412162 424102
rect 412218 424046 442758 424102
rect 442814 424046 442882 424102
rect 442938 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 499878 424102
rect 499934 424046 500002 424102
rect 500058 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 79878 423978
rect 79934 423922 80002 423978
rect 80058 423922 110598 423978
rect 110654 423922 110722 423978
rect 110778 423922 141318 423978
rect 141374 423922 141442 423978
rect 141498 423922 172038 423978
rect 172094 423922 172162 423978
rect 172218 423922 202758 423978
rect 202814 423922 202882 423978
rect 202938 423922 233478 423978
rect 233534 423922 233602 423978
rect 233658 423922 264198 423978
rect 264254 423922 264322 423978
rect 264378 423922 285714 423978
rect 285770 423922 285838 423978
rect 285894 423922 285962 423978
rect 286018 423922 286086 423978
rect 286142 423922 319878 423978
rect 319934 423922 320002 423978
rect 320058 423922 350598 423978
rect 350654 423922 350722 423978
rect 350778 423922 381318 423978
rect 381374 423922 381442 423978
rect 381498 423922 412038 423978
rect 412094 423922 412162 423978
rect 412218 423922 442758 423978
rect 442814 423922 442882 423978
rect 442938 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 499878 423978
rect 499934 423922 500002 423978
rect 500058 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect 56796 423478 283124 423494
rect 56796 423422 56812 423478
rect 56868 423422 283052 423478
rect 283108 423422 283124 423478
rect 56796 423406 283124 423422
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 64518 418350
rect 64574 418294 64642 418350
rect 64698 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 95238 418350
rect 95294 418294 95362 418350
rect 95418 418294 125958 418350
rect 126014 418294 126082 418350
rect 126138 418294 156678 418350
rect 156734 418294 156802 418350
rect 156858 418294 187398 418350
rect 187454 418294 187522 418350
rect 187578 418294 218118 418350
rect 218174 418294 218242 418350
rect 218298 418294 248838 418350
rect 248894 418294 248962 418350
rect 249018 418294 281994 418350
rect 282050 418294 282118 418350
rect 282174 418294 282242 418350
rect 282298 418294 282366 418350
rect 282422 418294 304518 418350
rect 304574 418294 304642 418350
rect 304698 418294 335238 418350
rect 335294 418294 335362 418350
rect 335418 418294 365958 418350
rect 366014 418294 366082 418350
rect 366138 418294 396678 418350
rect 396734 418294 396802 418350
rect 396858 418294 427398 418350
rect 427454 418294 427522 418350
rect 427578 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 484518 418350
rect 484574 418294 484642 418350
rect 484698 418294 515238 418350
rect 515294 418294 515362 418350
rect 515418 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 64518 418226
rect 64574 418170 64642 418226
rect 64698 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 95238 418226
rect 95294 418170 95362 418226
rect 95418 418170 125958 418226
rect 126014 418170 126082 418226
rect 126138 418170 156678 418226
rect 156734 418170 156802 418226
rect 156858 418170 187398 418226
rect 187454 418170 187522 418226
rect 187578 418170 218118 418226
rect 218174 418170 218242 418226
rect 218298 418170 248838 418226
rect 248894 418170 248962 418226
rect 249018 418170 281994 418226
rect 282050 418170 282118 418226
rect 282174 418170 282242 418226
rect 282298 418170 282366 418226
rect 282422 418170 304518 418226
rect 304574 418170 304642 418226
rect 304698 418170 335238 418226
rect 335294 418170 335362 418226
rect 335418 418170 365958 418226
rect 366014 418170 366082 418226
rect 366138 418170 396678 418226
rect 396734 418170 396802 418226
rect 396858 418170 427398 418226
rect 427454 418170 427522 418226
rect 427578 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 484518 418226
rect 484574 418170 484642 418226
rect 484698 418170 515238 418226
rect 515294 418170 515362 418226
rect 515418 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 64518 418102
rect 64574 418046 64642 418102
rect 64698 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 95238 418102
rect 95294 418046 95362 418102
rect 95418 418046 125958 418102
rect 126014 418046 126082 418102
rect 126138 418046 156678 418102
rect 156734 418046 156802 418102
rect 156858 418046 187398 418102
rect 187454 418046 187522 418102
rect 187578 418046 218118 418102
rect 218174 418046 218242 418102
rect 218298 418046 248838 418102
rect 248894 418046 248962 418102
rect 249018 418046 281994 418102
rect 282050 418046 282118 418102
rect 282174 418046 282242 418102
rect 282298 418046 282366 418102
rect 282422 418046 304518 418102
rect 304574 418046 304642 418102
rect 304698 418046 335238 418102
rect 335294 418046 335362 418102
rect 335418 418046 365958 418102
rect 366014 418046 366082 418102
rect 366138 418046 396678 418102
rect 396734 418046 396802 418102
rect 396858 418046 427398 418102
rect 427454 418046 427522 418102
rect 427578 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 484518 418102
rect 484574 418046 484642 418102
rect 484698 418046 515238 418102
rect 515294 418046 515362 418102
rect 515418 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 64518 417978
rect 64574 417922 64642 417978
rect 64698 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 95238 417978
rect 95294 417922 95362 417978
rect 95418 417922 125958 417978
rect 126014 417922 126082 417978
rect 126138 417922 156678 417978
rect 156734 417922 156802 417978
rect 156858 417922 187398 417978
rect 187454 417922 187522 417978
rect 187578 417922 218118 417978
rect 218174 417922 218242 417978
rect 218298 417922 248838 417978
rect 248894 417922 248962 417978
rect 249018 417922 281994 417978
rect 282050 417922 282118 417978
rect 282174 417922 282242 417978
rect 282298 417922 282366 417978
rect 282422 417922 304518 417978
rect 304574 417922 304642 417978
rect 304698 417922 335238 417978
rect 335294 417922 335362 417978
rect 335418 417922 365958 417978
rect 366014 417922 366082 417978
rect 366138 417922 396678 417978
rect 396734 417922 396802 417978
rect 396858 417922 427398 417978
rect 427454 417922 427522 417978
rect 427578 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 484518 417978
rect 484574 417922 484642 417978
rect 484698 417922 515238 417978
rect 515294 417922 515362 417978
rect 515418 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect 60156 409798 83652 409814
rect 60156 409742 60172 409798
rect 60228 409742 83580 409798
rect 83636 409742 83652 409798
rect 60156 409726 83652 409742
rect 60268 408178 83428 408194
rect 60268 408122 60284 408178
rect 60340 408122 83356 408178
rect 83412 408122 83428 408178
rect 60268 408106 83428 408122
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 79878 406350
rect 79934 406294 80002 406350
rect 80058 406294 110598 406350
rect 110654 406294 110722 406350
rect 110778 406294 141318 406350
rect 141374 406294 141442 406350
rect 141498 406294 172038 406350
rect 172094 406294 172162 406350
rect 172218 406294 202758 406350
rect 202814 406294 202882 406350
rect 202938 406294 233478 406350
rect 233534 406294 233602 406350
rect 233658 406294 264198 406350
rect 264254 406294 264322 406350
rect 264378 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 319878 406350
rect 319934 406294 320002 406350
rect 320058 406294 350598 406350
rect 350654 406294 350722 406350
rect 350778 406294 381318 406350
rect 381374 406294 381442 406350
rect 381498 406294 412038 406350
rect 412094 406294 412162 406350
rect 412218 406294 442758 406350
rect 442814 406294 442882 406350
rect 442938 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 499878 406350
rect 499934 406294 500002 406350
rect 500058 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 79878 406226
rect 79934 406170 80002 406226
rect 80058 406170 110598 406226
rect 110654 406170 110722 406226
rect 110778 406170 141318 406226
rect 141374 406170 141442 406226
rect 141498 406170 172038 406226
rect 172094 406170 172162 406226
rect 172218 406170 202758 406226
rect 202814 406170 202882 406226
rect 202938 406170 233478 406226
rect 233534 406170 233602 406226
rect 233658 406170 264198 406226
rect 264254 406170 264322 406226
rect 264378 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 319878 406226
rect 319934 406170 320002 406226
rect 320058 406170 350598 406226
rect 350654 406170 350722 406226
rect 350778 406170 381318 406226
rect 381374 406170 381442 406226
rect 381498 406170 412038 406226
rect 412094 406170 412162 406226
rect 412218 406170 442758 406226
rect 442814 406170 442882 406226
rect 442938 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 499878 406226
rect 499934 406170 500002 406226
rect 500058 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 79878 406102
rect 79934 406046 80002 406102
rect 80058 406046 110598 406102
rect 110654 406046 110722 406102
rect 110778 406046 141318 406102
rect 141374 406046 141442 406102
rect 141498 406046 172038 406102
rect 172094 406046 172162 406102
rect 172218 406046 202758 406102
rect 202814 406046 202882 406102
rect 202938 406046 233478 406102
rect 233534 406046 233602 406102
rect 233658 406046 264198 406102
rect 264254 406046 264322 406102
rect 264378 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 319878 406102
rect 319934 406046 320002 406102
rect 320058 406046 350598 406102
rect 350654 406046 350722 406102
rect 350778 406046 381318 406102
rect 381374 406046 381442 406102
rect 381498 406046 412038 406102
rect 412094 406046 412162 406102
rect 412218 406046 442758 406102
rect 442814 406046 442882 406102
rect 442938 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 499878 406102
rect 499934 406046 500002 406102
rect 500058 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 79878 405978
rect 79934 405922 80002 405978
rect 80058 405922 110598 405978
rect 110654 405922 110722 405978
rect 110778 405922 141318 405978
rect 141374 405922 141442 405978
rect 141498 405922 172038 405978
rect 172094 405922 172162 405978
rect 172218 405922 202758 405978
rect 202814 405922 202882 405978
rect 202938 405922 233478 405978
rect 233534 405922 233602 405978
rect 233658 405922 264198 405978
rect 264254 405922 264322 405978
rect 264378 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 319878 405978
rect 319934 405922 320002 405978
rect 320058 405922 350598 405978
rect 350654 405922 350722 405978
rect 350778 405922 381318 405978
rect 381374 405922 381442 405978
rect 381498 405922 412038 405978
rect 412094 405922 412162 405978
rect 412218 405922 442758 405978
rect 442814 405922 442882 405978
rect 442938 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 499878 405978
rect 499934 405922 500002 405978
rect 500058 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect 480604 405478 481700 405494
rect 480604 405422 480620 405478
rect 480676 405422 481628 405478
rect 481684 405422 481700 405478
rect 480604 405406 481700 405422
rect 60492 404758 83204 404774
rect 60492 404702 60508 404758
rect 60564 404702 83132 404758
rect 83188 404702 83204 404758
rect 60492 404686 83204 404702
rect 298604 404578 478564 404594
rect 298604 404522 298620 404578
rect 298676 404522 478492 404578
rect 478548 404522 478564 404578
rect 298604 404506 478564 404522
rect 303196 404398 468708 404414
rect 303196 404342 303212 404398
rect 303268 404342 467852 404398
rect 467908 404342 468636 404398
rect 468692 404342 468708 404398
rect 303196 404326 468708 404342
rect 260300 403138 481588 403154
rect 260300 403082 260316 403138
rect 260372 403082 481516 403138
rect 481572 403082 481588 403138
rect 260300 403066 481588 403082
rect 263660 402958 481476 402974
rect 263660 402902 263676 402958
rect 263732 402902 481404 402958
rect 481460 402902 481476 402958
rect 263660 402886 481476 402902
rect 298380 402778 483156 402794
rect 298380 402722 298396 402778
rect 298452 402722 483084 402778
rect 483140 402722 483156 402778
rect 298380 402706 483156 402722
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 64518 400350
rect 64574 400294 64642 400350
rect 64698 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 95238 400350
rect 95294 400294 95362 400350
rect 95418 400294 125958 400350
rect 126014 400294 126082 400350
rect 126138 400294 156678 400350
rect 156734 400294 156802 400350
rect 156858 400294 187398 400350
rect 187454 400294 187522 400350
rect 187578 400294 218118 400350
rect 218174 400294 218242 400350
rect 218298 400294 248838 400350
rect 248894 400294 248962 400350
rect 249018 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 374154 400350
rect 374210 400294 374278 400350
rect 374334 400294 374402 400350
rect 374458 400294 374526 400350
rect 374582 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 484518 400350
rect 484574 400294 484642 400350
rect 484698 400294 515238 400350
rect 515294 400294 515362 400350
rect 515418 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 64518 400226
rect 64574 400170 64642 400226
rect 64698 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 95238 400226
rect 95294 400170 95362 400226
rect 95418 400170 125958 400226
rect 126014 400170 126082 400226
rect 126138 400170 156678 400226
rect 156734 400170 156802 400226
rect 156858 400170 187398 400226
rect 187454 400170 187522 400226
rect 187578 400170 218118 400226
rect 218174 400170 218242 400226
rect 218298 400170 248838 400226
rect 248894 400170 248962 400226
rect 249018 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 374154 400226
rect 374210 400170 374278 400226
rect 374334 400170 374402 400226
rect 374458 400170 374526 400226
rect 374582 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 484518 400226
rect 484574 400170 484642 400226
rect 484698 400170 515238 400226
rect 515294 400170 515362 400226
rect 515418 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 64518 400102
rect 64574 400046 64642 400102
rect 64698 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 95238 400102
rect 95294 400046 95362 400102
rect 95418 400046 125958 400102
rect 126014 400046 126082 400102
rect 126138 400046 156678 400102
rect 156734 400046 156802 400102
rect 156858 400046 187398 400102
rect 187454 400046 187522 400102
rect 187578 400046 218118 400102
rect 218174 400046 218242 400102
rect 218298 400046 248838 400102
rect 248894 400046 248962 400102
rect 249018 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 374154 400102
rect 374210 400046 374278 400102
rect 374334 400046 374402 400102
rect 374458 400046 374526 400102
rect 374582 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 484518 400102
rect 484574 400046 484642 400102
rect 484698 400046 515238 400102
rect 515294 400046 515362 400102
rect 515418 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 64518 399978
rect 64574 399922 64642 399978
rect 64698 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 95238 399978
rect 95294 399922 95362 399978
rect 95418 399922 125958 399978
rect 126014 399922 126082 399978
rect 126138 399922 156678 399978
rect 156734 399922 156802 399978
rect 156858 399922 187398 399978
rect 187454 399922 187522 399978
rect 187578 399922 218118 399978
rect 218174 399922 218242 399978
rect 218298 399922 248838 399978
rect 248894 399922 248962 399978
rect 249018 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 374154 399978
rect 374210 399922 374278 399978
rect 374334 399922 374402 399978
rect 374458 399922 374526 399978
rect 374582 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 484518 399978
rect 484574 399922 484642 399978
rect 484698 399922 515238 399978
rect 515294 399922 515362 399978
rect 515418 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect 298716 398098 483044 398114
rect 298716 398042 298732 398098
rect 298788 398042 482972 398098
rect 483028 398042 483044 398098
rect 298716 398026 483044 398042
rect 273516 388918 526724 388934
rect 273516 388862 273532 388918
rect 273588 388862 525868 388918
rect 525924 388862 526652 388918
rect 526708 388862 526724 388918
rect 273516 388846 526724 388862
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 79878 388350
rect 79934 388294 80002 388350
rect 80058 388294 110598 388350
rect 110654 388294 110722 388350
rect 110778 388294 141318 388350
rect 141374 388294 141442 388350
rect 141498 388294 172038 388350
rect 172094 388294 172162 388350
rect 172218 388294 202758 388350
rect 202814 388294 202882 388350
rect 202938 388294 233478 388350
rect 233534 388294 233602 388350
rect 233658 388294 264198 388350
rect 264254 388294 264322 388350
rect 264378 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 377874 388350
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388294 499878 388350
rect 499934 388294 500002 388350
rect 500058 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 79878 388226
rect 79934 388170 80002 388226
rect 80058 388170 110598 388226
rect 110654 388170 110722 388226
rect 110778 388170 141318 388226
rect 141374 388170 141442 388226
rect 141498 388170 172038 388226
rect 172094 388170 172162 388226
rect 172218 388170 202758 388226
rect 202814 388170 202882 388226
rect 202938 388170 233478 388226
rect 233534 388170 233602 388226
rect 233658 388170 264198 388226
rect 264254 388170 264322 388226
rect 264378 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 499878 388226
rect 499934 388170 500002 388226
rect 500058 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 79878 388102
rect 79934 388046 80002 388102
rect 80058 388046 110598 388102
rect 110654 388046 110722 388102
rect 110778 388046 141318 388102
rect 141374 388046 141442 388102
rect 141498 388046 172038 388102
rect 172094 388046 172162 388102
rect 172218 388046 202758 388102
rect 202814 388046 202882 388102
rect 202938 388046 233478 388102
rect 233534 388046 233602 388102
rect 233658 388046 264198 388102
rect 264254 388046 264322 388102
rect 264378 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 499878 388102
rect 499934 388046 500002 388102
rect 500058 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 79878 387978
rect 79934 387922 80002 387978
rect 80058 387922 110598 387978
rect 110654 387922 110722 387978
rect 110778 387922 141318 387978
rect 141374 387922 141442 387978
rect 141498 387922 172038 387978
rect 172094 387922 172162 387978
rect 172218 387922 202758 387978
rect 202814 387922 202882 387978
rect 202938 387922 233478 387978
rect 233534 387922 233602 387978
rect 233658 387922 264198 387978
rect 264254 387922 264322 387978
rect 264378 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 499878 387978
rect 499934 387922 500002 387978
rect 500058 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect 276428 387658 591124 387674
rect 276428 387602 276444 387658
rect 276500 387602 591052 387658
rect 591108 387602 591124 387658
rect 276428 387586 591124 387602
rect 60268 383158 84884 383174
rect 60268 383102 60284 383158
rect 60340 383102 84812 383158
rect 84868 383102 84884 383158
rect 60268 383086 84884 383102
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 64518 382350
rect 64574 382294 64642 382350
rect 64698 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 95238 382350
rect 95294 382294 95362 382350
rect 95418 382294 125958 382350
rect 126014 382294 126082 382350
rect 126138 382294 156678 382350
rect 156734 382294 156802 382350
rect 156858 382294 187398 382350
rect 187454 382294 187522 382350
rect 187578 382294 218118 382350
rect 218174 382294 218242 382350
rect 218298 382294 248838 382350
rect 248894 382294 248962 382350
rect 249018 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 374154 382350
rect 374210 382294 374278 382350
rect 374334 382294 374402 382350
rect 374458 382294 374526 382350
rect 374582 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 64518 382226
rect 64574 382170 64642 382226
rect 64698 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 95238 382226
rect 95294 382170 95362 382226
rect 95418 382170 125958 382226
rect 126014 382170 126082 382226
rect 126138 382170 156678 382226
rect 156734 382170 156802 382226
rect 156858 382170 187398 382226
rect 187454 382170 187522 382226
rect 187578 382170 218118 382226
rect 218174 382170 218242 382226
rect 218298 382170 248838 382226
rect 248894 382170 248962 382226
rect 249018 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 374154 382226
rect 374210 382170 374278 382226
rect 374334 382170 374402 382226
rect 374458 382170 374526 382226
rect 374582 382170 404874 382226
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 64518 382102
rect 64574 382046 64642 382102
rect 64698 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 95238 382102
rect 95294 382046 95362 382102
rect 95418 382046 125958 382102
rect 126014 382046 126082 382102
rect 126138 382046 156678 382102
rect 156734 382046 156802 382102
rect 156858 382046 187398 382102
rect 187454 382046 187522 382102
rect 187578 382046 218118 382102
rect 218174 382046 218242 382102
rect 218298 382046 248838 382102
rect 248894 382046 248962 382102
rect 249018 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 374154 382102
rect 374210 382046 374278 382102
rect 374334 382046 374402 382102
rect 374458 382046 374526 382102
rect 374582 382046 404874 382102
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 64518 381978
rect 64574 381922 64642 381978
rect 64698 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 95238 381978
rect 95294 381922 95362 381978
rect 95418 381922 125958 381978
rect 126014 381922 126082 381978
rect 126138 381922 156678 381978
rect 156734 381922 156802 381978
rect 156858 381922 187398 381978
rect 187454 381922 187522 381978
rect 187578 381922 218118 381978
rect 218174 381922 218242 381978
rect 218298 381922 248838 381978
rect 248894 381922 248962 381978
rect 249018 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 374154 381978
rect 374210 381922 374278 381978
rect 374334 381922 374402 381978
rect 374458 381922 374526 381978
rect 374582 381922 404874 381978
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect 289868 377938 521124 377954
rect 289868 377882 289884 377938
rect 289940 377882 521052 377938
rect 521108 377882 521124 377938
rect 289868 377866 521124 377882
rect 293116 377758 494916 377774
rect 293116 377702 293132 377758
rect 293188 377702 494844 377758
rect 494900 377702 494916 377758
rect 293116 377686 494916 377702
rect 296588 377578 498948 377594
rect 296588 377522 296604 377578
rect 296660 377522 498876 377578
rect 498932 377522 498948 377578
rect 296588 377506 498948 377522
rect 278220 376498 590228 376514
rect 278220 376442 278236 376498
rect 278292 376442 590156 376498
rect 590212 376442 590228 376498
rect 278220 376426 590228 376442
rect 60716 374878 83204 374894
rect 60716 374822 60732 374878
rect 60788 374822 83132 374878
rect 83188 374822 83204 374878
rect 60716 374806 83204 374822
rect 60156 374698 83428 374714
rect 60156 374642 60172 374698
rect 60228 374642 83356 374698
rect 83412 374642 83428 374698
rect 60156 374626 83428 374642
rect 295244 373798 505780 373814
rect 295244 373742 295260 373798
rect 295316 373742 505708 373798
rect 505764 373742 505780 373798
rect 295244 373726 505780 373742
rect 273740 371458 451236 371474
rect 273740 371402 273756 371458
rect 273812 371402 451164 371458
rect 451220 371402 451236 371458
rect 273740 371386 451236 371402
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 79878 370350
rect 79934 370294 80002 370350
rect 80058 370294 110598 370350
rect 110654 370294 110722 370350
rect 110778 370294 141318 370350
rect 141374 370294 141442 370350
rect 141498 370294 172038 370350
rect 172094 370294 172162 370350
rect 172218 370294 202758 370350
rect 202814 370294 202882 370350
rect 202938 370294 233478 370350
rect 233534 370294 233602 370350
rect 233658 370294 264198 370350
rect 264254 370294 264322 370350
rect 264378 370294 285714 370350
rect 285770 370294 285838 370350
rect 285894 370294 285962 370350
rect 286018 370294 286086 370350
rect 286142 370294 301932 370350
rect 301988 370294 302056 370350
rect 302112 370294 302180 370350
rect 302236 370294 302304 370350
rect 302360 370294 316434 370350
rect 316490 370294 316558 370350
rect 316614 370294 316682 370350
rect 316738 370294 316806 370350
rect 316862 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 386614 370350
rect 386670 370294 386738 370350
rect 386794 370294 386862 370350
rect 386918 370294 386986 370350
rect 387042 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 79878 370226
rect 79934 370170 80002 370226
rect 80058 370170 110598 370226
rect 110654 370170 110722 370226
rect 110778 370170 141318 370226
rect 141374 370170 141442 370226
rect 141498 370170 172038 370226
rect 172094 370170 172162 370226
rect 172218 370170 202758 370226
rect 202814 370170 202882 370226
rect 202938 370170 233478 370226
rect 233534 370170 233602 370226
rect 233658 370170 264198 370226
rect 264254 370170 264322 370226
rect 264378 370170 285714 370226
rect 285770 370170 285838 370226
rect 285894 370170 285962 370226
rect 286018 370170 286086 370226
rect 286142 370170 301932 370226
rect 301988 370170 302056 370226
rect 302112 370170 302180 370226
rect 302236 370170 302304 370226
rect 302360 370170 316434 370226
rect 316490 370170 316558 370226
rect 316614 370170 316682 370226
rect 316738 370170 316806 370226
rect 316862 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 386614 370226
rect 386670 370170 386738 370226
rect 386794 370170 386862 370226
rect 386918 370170 386986 370226
rect 387042 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 79878 370102
rect 79934 370046 80002 370102
rect 80058 370046 110598 370102
rect 110654 370046 110722 370102
rect 110778 370046 141318 370102
rect 141374 370046 141442 370102
rect 141498 370046 172038 370102
rect 172094 370046 172162 370102
rect 172218 370046 202758 370102
rect 202814 370046 202882 370102
rect 202938 370046 233478 370102
rect 233534 370046 233602 370102
rect 233658 370046 264198 370102
rect 264254 370046 264322 370102
rect 264378 370046 285714 370102
rect 285770 370046 285838 370102
rect 285894 370046 285962 370102
rect 286018 370046 286086 370102
rect 286142 370046 301932 370102
rect 301988 370046 302056 370102
rect 302112 370046 302180 370102
rect 302236 370046 302304 370102
rect 302360 370046 316434 370102
rect 316490 370046 316558 370102
rect 316614 370046 316682 370102
rect 316738 370046 316806 370102
rect 316862 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 386614 370102
rect 386670 370046 386738 370102
rect 386794 370046 386862 370102
rect 386918 370046 386986 370102
rect 387042 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 79878 369978
rect 79934 369922 80002 369978
rect 80058 369922 110598 369978
rect 110654 369922 110722 369978
rect 110778 369922 141318 369978
rect 141374 369922 141442 369978
rect 141498 369922 172038 369978
rect 172094 369922 172162 369978
rect 172218 369922 202758 369978
rect 202814 369922 202882 369978
rect 202938 369922 233478 369978
rect 233534 369922 233602 369978
rect 233658 369922 264198 369978
rect 264254 369922 264322 369978
rect 264378 369922 285714 369978
rect 285770 369922 285838 369978
rect 285894 369922 285962 369978
rect 286018 369922 286086 369978
rect 286142 369922 301932 369978
rect 301988 369922 302056 369978
rect 302112 369922 302180 369978
rect 302236 369922 302304 369978
rect 302360 369922 316434 369978
rect 316490 369922 316558 369978
rect 316614 369922 316682 369978
rect 316738 369922 316806 369978
rect 316862 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 386614 369978
rect 386670 369922 386738 369978
rect 386794 369922 386862 369978
rect 386918 369922 386986 369978
rect 387042 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect 295020 368758 502420 368774
rect 295020 368702 295036 368758
rect 295092 368702 502348 368758
rect 502404 368702 502420 368758
rect 295020 368686 502420 368702
rect 60156 368218 83652 368234
rect 60156 368162 60172 368218
rect 60228 368162 83580 368218
rect 83636 368162 83652 368218
rect 60156 368146 83652 368162
rect 60716 368038 83876 368054
rect 60716 367982 60732 368038
rect 60788 367982 83804 368038
rect 83860 367982 83876 368038
rect 60716 367966 83876 367982
rect 273740 368038 457956 368054
rect 273740 367982 273756 368038
rect 273812 367982 457884 368038
rect 457940 367982 457956 368038
rect 273740 367966 457956 367982
rect 60716 366418 83764 366434
rect 60716 366362 60732 366418
rect 60788 366362 83692 366418
rect 83748 366362 83764 366418
rect 60716 366346 83764 366362
rect 273740 366418 454596 366434
rect 273740 366362 273756 366418
rect 273812 366362 454524 366418
rect 454580 366362 454596 366418
rect 273740 366346 454596 366362
rect 273740 364798 451124 364814
rect 273740 364742 273756 364798
rect 273812 364742 451052 364798
rect 451108 364742 451124 364798
rect 273740 364726 451124 364742
rect 273740 364618 454484 364634
rect 273740 364562 273756 364618
rect 273812 364562 454412 364618
rect 454468 364562 454484 364618
rect 273740 364546 454484 364562
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 64518 364350
rect 64574 364294 64642 364350
rect 64698 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 95238 364350
rect 95294 364294 95362 364350
rect 95418 364294 125958 364350
rect 126014 364294 126082 364350
rect 126138 364294 156678 364350
rect 156734 364294 156802 364350
rect 156858 364294 187398 364350
rect 187454 364294 187522 364350
rect 187578 364294 218118 364350
rect 218174 364294 218242 364350
rect 218298 364294 248838 364350
rect 248894 364294 248962 364350
rect 249018 364294 281994 364350
rect 282050 364294 282118 364350
rect 282174 364294 282242 364350
rect 282298 364294 282366 364350
rect 282422 364294 302732 364350
rect 302788 364294 302856 364350
rect 302912 364294 302980 364350
rect 303036 364294 303104 364350
rect 303160 364294 312714 364350
rect 312770 364294 312838 364350
rect 312894 364294 312962 364350
rect 313018 364294 313086 364350
rect 313142 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 374154 364350
rect 374210 364294 374278 364350
rect 374334 364294 374402 364350
rect 374458 364294 374526 364350
rect 374582 364294 387414 364350
rect 387470 364294 387538 364350
rect 387594 364294 387662 364350
rect 387718 364294 387786 364350
rect 387842 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 64518 364226
rect 64574 364170 64642 364226
rect 64698 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 95238 364226
rect 95294 364170 95362 364226
rect 95418 364170 125958 364226
rect 126014 364170 126082 364226
rect 126138 364170 156678 364226
rect 156734 364170 156802 364226
rect 156858 364170 187398 364226
rect 187454 364170 187522 364226
rect 187578 364170 218118 364226
rect 218174 364170 218242 364226
rect 218298 364170 248838 364226
rect 248894 364170 248962 364226
rect 249018 364170 281994 364226
rect 282050 364170 282118 364226
rect 282174 364170 282242 364226
rect 282298 364170 282366 364226
rect 282422 364170 302732 364226
rect 302788 364170 302856 364226
rect 302912 364170 302980 364226
rect 303036 364170 303104 364226
rect 303160 364170 312714 364226
rect 312770 364170 312838 364226
rect 312894 364170 312962 364226
rect 313018 364170 313086 364226
rect 313142 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 374154 364226
rect 374210 364170 374278 364226
rect 374334 364170 374402 364226
rect 374458 364170 374526 364226
rect 374582 364170 387414 364226
rect 387470 364170 387538 364226
rect 387594 364170 387662 364226
rect 387718 364170 387786 364226
rect 387842 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 64518 364102
rect 64574 364046 64642 364102
rect 64698 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 95238 364102
rect 95294 364046 95362 364102
rect 95418 364046 125958 364102
rect 126014 364046 126082 364102
rect 126138 364046 156678 364102
rect 156734 364046 156802 364102
rect 156858 364046 187398 364102
rect 187454 364046 187522 364102
rect 187578 364046 218118 364102
rect 218174 364046 218242 364102
rect 218298 364046 248838 364102
rect 248894 364046 248962 364102
rect 249018 364046 281994 364102
rect 282050 364046 282118 364102
rect 282174 364046 282242 364102
rect 282298 364046 282366 364102
rect 282422 364046 302732 364102
rect 302788 364046 302856 364102
rect 302912 364046 302980 364102
rect 303036 364046 303104 364102
rect 303160 364046 312714 364102
rect 312770 364046 312838 364102
rect 312894 364046 312962 364102
rect 313018 364046 313086 364102
rect 313142 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 374154 364102
rect 374210 364046 374278 364102
rect 374334 364046 374402 364102
rect 374458 364046 374526 364102
rect 374582 364046 387414 364102
rect 387470 364046 387538 364102
rect 387594 364046 387662 364102
rect 387718 364046 387786 364102
rect 387842 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 64518 363978
rect 64574 363922 64642 363978
rect 64698 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 95238 363978
rect 95294 363922 95362 363978
rect 95418 363922 125958 363978
rect 126014 363922 126082 363978
rect 126138 363922 156678 363978
rect 156734 363922 156802 363978
rect 156858 363922 187398 363978
rect 187454 363922 187522 363978
rect 187578 363922 218118 363978
rect 218174 363922 218242 363978
rect 218298 363922 248838 363978
rect 248894 363922 248962 363978
rect 249018 363922 281994 363978
rect 282050 363922 282118 363978
rect 282174 363922 282242 363978
rect 282298 363922 282366 363978
rect 282422 363922 302732 363978
rect 302788 363922 302856 363978
rect 302912 363922 302980 363978
rect 303036 363922 303104 363978
rect 303160 363922 312714 363978
rect 312770 363922 312838 363978
rect 312894 363922 312962 363978
rect 313018 363922 313086 363978
rect 313142 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 374154 363978
rect 374210 363922 374278 363978
rect 374334 363922 374402 363978
rect 374458 363922 374526 363978
rect 374582 363922 387414 363978
rect 387470 363922 387538 363978
rect 387594 363922 387662 363978
rect 387718 363922 387786 363978
rect 387842 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect 273740 361378 456276 361394
rect 273740 361322 273756 361378
rect 273812 361322 456204 361378
rect 456260 361322 456276 361378
rect 273740 361306 456276 361322
rect 294908 360298 499060 360314
rect 294908 360242 294924 360298
rect 294980 360242 498988 360298
rect 499044 360242 499060 360298
rect 294908 360226 499060 360242
rect 273740 358678 452804 358694
rect 273740 358622 273756 358678
rect 273812 358622 452732 358678
rect 452788 358622 452804 358678
rect 273740 358606 452804 358622
rect 273740 356338 452916 356354
rect 273740 356282 273756 356338
rect 273812 356282 452844 356338
rect 452900 356282 452916 356338
rect 273740 356266 452916 356282
rect 273740 354538 449556 354554
rect 273740 354482 273756 354538
rect 273812 354482 449484 354538
rect 449540 354482 449556 354538
rect 273740 354466 449556 354482
rect 273740 353638 456164 353654
rect 273740 353582 273756 353638
rect 273812 353582 456092 353638
rect 456148 353582 456164 353638
rect 273740 353566 456164 353582
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 79878 352350
rect 79934 352294 80002 352350
rect 80058 352294 110598 352350
rect 110654 352294 110722 352350
rect 110778 352294 141318 352350
rect 141374 352294 141442 352350
rect 141498 352294 172038 352350
rect 172094 352294 172162 352350
rect 172218 352294 202758 352350
rect 202814 352294 202882 352350
rect 202938 352294 233478 352350
rect 233534 352294 233602 352350
rect 233658 352294 264198 352350
rect 264254 352294 264322 352350
rect 264378 352294 285714 352350
rect 285770 352294 285838 352350
rect 285894 352294 285962 352350
rect 286018 352294 286086 352350
rect 286142 352294 301932 352350
rect 301988 352294 302056 352350
rect 302112 352294 302180 352350
rect 302236 352294 302304 352350
rect 302360 352294 316434 352350
rect 316490 352294 316558 352350
rect 316614 352294 316682 352350
rect 316738 352294 316806 352350
rect 316862 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 386614 352350
rect 386670 352294 386738 352350
rect 386794 352294 386862 352350
rect 386918 352294 386986 352350
rect 387042 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 79878 352226
rect 79934 352170 80002 352226
rect 80058 352170 110598 352226
rect 110654 352170 110722 352226
rect 110778 352170 141318 352226
rect 141374 352170 141442 352226
rect 141498 352170 172038 352226
rect 172094 352170 172162 352226
rect 172218 352170 202758 352226
rect 202814 352170 202882 352226
rect 202938 352170 233478 352226
rect 233534 352170 233602 352226
rect 233658 352170 264198 352226
rect 264254 352170 264322 352226
rect 264378 352170 285714 352226
rect 285770 352170 285838 352226
rect 285894 352170 285962 352226
rect 286018 352170 286086 352226
rect 286142 352170 301932 352226
rect 301988 352170 302056 352226
rect 302112 352170 302180 352226
rect 302236 352170 302304 352226
rect 302360 352170 316434 352226
rect 316490 352170 316558 352226
rect 316614 352170 316682 352226
rect 316738 352170 316806 352226
rect 316862 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 386614 352226
rect 386670 352170 386738 352226
rect 386794 352170 386862 352226
rect 386918 352170 386986 352226
rect 387042 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 79878 352102
rect 79934 352046 80002 352102
rect 80058 352046 110598 352102
rect 110654 352046 110722 352102
rect 110778 352046 141318 352102
rect 141374 352046 141442 352102
rect 141498 352046 172038 352102
rect 172094 352046 172162 352102
rect 172218 352046 202758 352102
rect 202814 352046 202882 352102
rect 202938 352046 233478 352102
rect 233534 352046 233602 352102
rect 233658 352046 264198 352102
rect 264254 352046 264322 352102
rect 264378 352046 285714 352102
rect 285770 352046 285838 352102
rect 285894 352046 285962 352102
rect 286018 352046 286086 352102
rect 286142 352046 301932 352102
rect 301988 352046 302056 352102
rect 302112 352046 302180 352102
rect 302236 352046 302304 352102
rect 302360 352046 316434 352102
rect 316490 352046 316558 352102
rect 316614 352046 316682 352102
rect 316738 352046 316806 352102
rect 316862 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 386614 352102
rect 386670 352046 386738 352102
rect 386794 352046 386862 352102
rect 386918 352046 386986 352102
rect 387042 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 79878 351978
rect 79934 351922 80002 351978
rect 80058 351922 110598 351978
rect 110654 351922 110722 351978
rect 110778 351922 141318 351978
rect 141374 351922 141442 351978
rect 141498 351922 172038 351978
rect 172094 351922 172162 351978
rect 172218 351922 202758 351978
rect 202814 351922 202882 351978
rect 202938 351922 233478 351978
rect 233534 351922 233602 351978
rect 233658 351922 264198 351978
rect 264254 351922 264322 351978
rect 264378 351922 285714 351978
rect 285770 351922 285838 351978
rect 285894 351922 285962 351978
rect 286018 351922 286086 351978
rect 286142 351922 301932 351978
rect 301988 351922 302056 351978
rect 302112 351922 302180 351978
rect 302236 351922 302304 351978
rect 302360 351922 316434 351978
rect 316490 351922 316558 351978
rect 316614 351922 316682 351978
rect 316738 351922 316806 351978
rect 316862 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 386614 351978
rect 386670 351922 386738 351978
rect 386794 351922 386862 351978
rect 386918 351922 386986 351978
rect 387042 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect 273292 350218 457844 350234
rect 273292 350162 273308 350218
rect 273364 350162 457772 350218
rect 457828 350162 457844 350218
rect 273292 350146 457844 350162
rect 60492 350038 69764 350054
rect 60492 349982 60508 350038
rect 60564 349982 69692 350038
rect 69748 349982 69764 350038
rect 60492 349966 69764 349982
rect 273740 349498 355364 349514
rect 273740 349442 273756 349498
rect 273812 349442 355292 349498
rect 355348 349442 355364 349498
rect 273740 349426 355364 349442
rect 294796 348598 496036 348614
rect 294796 348542 294812 348598
rect 294868 348542 495964 348598
rect 496020 348542 496036 348598
rect 294796 348526 496036 348542
rect 4156 347698 83540 347714
rect 4156 347642 4172 347698
rect 4228 347642 83468 347698
rect 83524 347642 83540 347698
rect 4156 347626 83540 347642
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 64518 346350
rect 64574 346294 64642 346350
rect 64698 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 95238 346350
rect 95294 346294 95362 346350
rect 95418 346294 125958 346350
rect 126014 346294 126082 346350
rect 126138 346294 156678 346350
rect 156734 346294 156802 346350
rect 156858 346294 187398 346350
rect 187454 346294 187522 346350
rect 187578 346294 218118 346350
rect 218174 346294 218242 346350
rect 218298 346294 248838 346350
rect 248894 346294 248962 346350
rect 249018 346294 281994 346350
rect 282050 346294 282118 346350
rect 282174 346294 282242 346350
rect 282298 346294 282366 346350
rect 282422 346294 302732 346350
rect 302788 346294 302856 346350
rect 302912 346294 302980 346350
rect 303036 346294 303104 346350
rect 303160 346294 312714 346350
rect 312770 346294 312838 346350
rect 312894 346294 312962 346350
rect 313018 346294 313086 346350
rect 313142 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 374154 346350
rect 374210 346294 374278 346350
rect 374334 346294 374402 346350
rect 374458 346294 374526 346350
rect 374582 346294 387414 346350
rect 387470 346294 387538 346350
rect 387594 346294 387662 346350
rect 387718 346294 387786 346350
rect 387842 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 64518 346226
rect 64574 346170 64642 346226
rect 64698 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 95238 346226
rect 95294 346170 95362 346226
rect 95418 346170 125958 346226
rect 126014 346170 126082 346226
rect 126138 346170 156678 346226
rect 156734 346170 156802 346226
rect 156858 346170 187398 346226
rect 187454 346170 187522 346226
rect 187578 346170 218118 346226
rect 218174 346170 218242 346226
rect 218298 346170 248838 346226
rect 248894 346170 248962 346226
rect 249018 346170 281994 346226
rect 282050 346170 282118 346226
rect 282174 346170 282242 346226
rect 282298 346170 282366 346226
rect 282422 346170 302732 346226
rect 302788 346170 302856 346226
rect 302912 346170 302980 346226
rect 303036 346170 303104 346226
rect 303160 346170 312714 346226
rect 312770 346170 312838 346226
rect 312894 346170 312962 346226
rect 313018 346170 313086 346226
rect 313142 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 374154 346226
rect 374210 346170 374278 346226
rect 374334 346170 374402 346226
rect 374458 346170 374526 346226
rect 374582 346170 387414 346226
rect 387470 346170 387538 346226
rect 387594 346170 387662 346226
rect 387718 346170 387786 346226
rect 387842 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 64518 346102
rect 64574 346046 64642 346102
rect 64698 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 95238 346102
rect 95294 346046 95362 346102
rect 95418 346046 125958 346102
rect 126014 346046 126082 346102
rect 126138 346046 156678 346102
rect 156734 346046 156802 346102
rect 156858 346046 187398 346102
rect 187454 346046 187522 346102
rect 187578 346046 218118 346102
rect 218174 346046 218242 346102
rect 218298 346046 248838 346102
rect 248894 346046 248962 346102
rect 249018 346046 281994 346102
rect 282050 346046 282118 346102
rect 282174 346046 282242 346102
rect 282298 346046 282366 346102
rect 282422 346046 302732 346102
rect 302788 346046 302856 346102
rect 302912 346046 302980 346102
rect 303036 346046 303104 346102
rect 303160 346046 312714 346102
rect 312770 346046 312838 346102
rect 312894 346046 312962 346102
rect 313018 346046 313086 346102
rect 313142 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 374154 346102
rect 374210 346046 374278 346102
rect 374334 346046 374402 346102
rect 374458 346046 374526 346102
rect 374582 346046 387414 346102
rect 387470 346046 387538 346102
rect 387594 346046 387662 346102
rect 387718 346046 387786 346102
rect 387842 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 64518 345978
rect 64574 345922 64642 345978
rect 64698 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 95238 345978
rect 95294 345922 95362 345978
rect 95418 345922 125958 345978
rect 126014 345922 126082 345978
rect 126138 345922 156678 345978
rect 156734 345922 156802 345978
rect 156858 345922 187398 345978
rect 187454 345922 187522 345978
rect 187578 345922 218118 345978
rect 218174 345922 218242 345978
rect 218298 345922 248838 345978
rect 248894 345922 248962 345978
rect 249018 345922 281994 345978
rect 282050 345922 282118 345978
rect 282174 345922 282242 345978
rect 282298 345922 282366 345978
rect 282422 345922 302732 345978
rect 302788 345922 302856 345978
rect 302912 345922 302980 345978
rect 303036 345922 303104 345978
rect 303160 345922 312714 345978
rect 312770 345922 312838 345978
rect 312894 345922 312962 345978
rect 313018 345922 313086 345978
rect 313142 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 374154 345978
rect 374210 345922 374278 345978
rect 374334 345922 374402 345978
rect 374458 345922 374526 345978
rect 374582 345922 387414 345978
rect 387470 345922 387538 345978
rect 387594 345922 387662 345978
rect 387718 345922 387786 345978
rect 387842 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect 281356 345718 519556 345734
rect 281356 345662 281372 345718
rect 281428 345662 519484 345718
rect 519540 345662 519556 345718
rect 281356 345646 519556 345662
rect 289756 345538 516196 345554
rect 289756 345482 289772 345538
rect 289828 345482 516124 345538
rect 516180 345482 516196 345538
rect 289756 345466 516196 345482
rect 284940 345358 509476 345374
rect 284940 345302 284956 345358
rect 285012 345302 509404 345358
rect 509460 345302 509476 345358
rect 284940 345286 509476 345302
rect 296476 345178 512836 345194
rect 296476 345122 296492 345178
rect 296548 345122 512764 345178
rect 512820 345122 512836 345178
rect 296476 345106 512836 345122
rect 60492 344458 78164 344474
rect 60492 344402 60508 344458
rect 60564 344402 78092 344458
rect 78148 344402 78164 344458
rect 60492 344386 78164 344402
rect 273740 343738 358724 343754
rect 273740 343682 273756 343738
rect 273812 343682 358652 343738
rect 358708 343682 358724 343738
rect 273740 343666 358724 343682
rect 273068 343558 449444 343574
rect 273068 343502 273084 343558
rect 273140 343502 449372 343558
rect 449428 343502 449444 343558
rect 273068 343486 449444 343502
rect 273628 341938 447540 341954
rect 273628 341882 273644 341938
rect 273700 341882 447468 341938
rect 447524 341882 447540 341938
rect 273628 341866 447540 341882
rect 301068 340318 475764 340334
rect 301068 340262 301084 340318
rect 301140 340262 475692 340318
rect 475748 340262 475764 340318
rect 301068 340246 475764 340262
rect 300844 340138 476324 340154
rect 300844 340082 300860 340138
rect 300916 340082 476252 340138
rect 476308 340082 476324 340138
rect 300844 340066 476324 340082
rect 288076 339238 475540 339254
rect 288076 339182 288092 339238
rect 288148 339182 475468 339238
rect 475524 339182 475540 339238
rect 288076 339166 475540 339182
rect 279676 337618 475540 337634
rect 279676 337562 279692 337618
rect 279748 337562 475468 337618
rect 475524 337562 475540 337618
rect 279676 337546 475540 337562
rect 298268 337438 475652 337454
rect 298268 337382 298284 337438
rect 298340 337382 475580 337438
rect 475636 337382 475652 337438
rect 298268 337366 475652 337382
rect 60156 335998 83316 336014
rect 60156 335942 60172 335998
rect 60228 335942 83244 335998
rect 83300 335942 83316 335998
rect 60156 335926 83316 335942
rect 278108 335998 475540 336014
rect 278108 335942 278124 335998
rect 278180 335942 475468 335998
rect 475524 335942 475540 335998
rect 278108 335926 475540 335942
rect 60716 335818 80292 335834
rect 60716 335762 60732 335818
rect 60788 335762 80220 335818
rect 80276 335762 80292 335818
rect 60716 335746 80292 335762
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 79878 334350
rect 79934 334294 80002 334350
rect 80058 334294 110598 334350
rect 110654 334294 110722 334350
rect 110778 334294 141318 334350
rect 141374 334294 141442 334350
rect 141498 334294 172038 334350
rect 172094 334294 172162 334350
rect 172218 334294 202758 334350
rect 202814 334294 202882 334350
rect 202938 334294 233478 334350
rect 233534 334294 233602 334350
rect 233658 334294 264198 334350
rect 264254 334294 264322 334350
rect 264378 334294 285714 334350
rect 285770 334294 285838 334350
rect 285894 334294 285962 334350
rect 286018 334294 286086 334350
rect 286142 334294 301932 334350
rect 301988 334294 302056 334350
rect 302112 334294 302180 334350
rect 302236 334294 302304 334350
rect 302360 334294 316434 334350
rect 316490 334294 316558 334350
rect 316614 334294 316682 334350
rect 316738 334294 316806 334350
rect 316862 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 386614 334350
rect 386670 334294 386738 334350
rect 386794 334294 386862 334350
rect 386918 334294 386986 334350
rect 387042 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 499878 334350
rect 499934 334294 500002 334350
rect 500058 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 79878 334226
rect 79934 334170 80002 334226
rect 80058 334170 110598 334226
rect 110654 334170 110722 334226
rect 110778 334170 141318 334226
rect 141374 334170 141442 334226
rect 141498 334170 172038 334226
rect 172094 334170 172162 334226
rect 172218 334170 202758 334226
rect 202814 334170 202882 334226
rect 202938 334170 233478 334226
rect 233534 334170 233602 334226
rect 233658 334170 264198 334226
rect 264254 334170 264322 334226
rect 264378 334170 285714 334226
rect 285770 334170 285838 334226
rect 285894 334170 285962 334226
rect 286018 334170 286086 334226
rect 286142 334170 301932 334226
rect 301988 334170 302056 334226
rect 302112 334170 302180 334226
rect 302236 334170 302304 334226
rect 302360 334170 316434 334226
rect 316490 334170 316558 334226
rect 316614 334170 316682 334226
rect 316738 334170 316806 334226
rect 316862 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 386614 334226
rect 386670 334170 386738 334226
rect 386794 334170 386862 334226
rect 386918 334170 386986 334226
rect 387042 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 499878 334226
rect 499934 334170 500002 334226
rect 500058 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 79878 334102
rect 79934 334046 80002 334102
rect 80058 334046 110598 334102
rect 110654 334046 110722 334102
rect 110778 334046 141318 334102
rect 141374 334046 141442 334102
rect 141498 334046 172038 334102
rect 172094 334046 172162 334102
rect 172218 334046 202758 334102
rect 202814 334046 202882 334102
rect 202938 334046 233478 334102
rect 233534 334046 233602 334102
rect 233658 334046 264198 334102
rect 264254 334046 264322 334102
rect 264378 334046 285714 334102
rect 285770 334046 285838 334102
rect 285894 334046 285962 334102
rect 286018 334046 286086 334102
rect 286142 334046 301932 334102
rect 301988 334046 302056 334102
rect 302112 334046 302180 334102
rect 302236 334046 302304 334102
rect 302360 334046 316434 334102
rect 316490 334046 316558 334102
rect 316614 334046 316682 334102
rect 316738 334046 316806 334102
rect 316862 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 386614 334102
rect 386670 334046 386738 334102
rect 386794 334046 386862 334102
rect 386918 334046 386986 334102
rect 387042 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 499878 334102
rect 499934 334046 500002 334102
rect 500058 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 79878 333978
rect 79934 333922 80002 333978
rect 80058 333922 110598 333978
rect 110654 333922 110722 333978
rect 110778 333922 141318 333978
rect 141374 333922 141442 333978
rect 141498 333922 172038 333978
rect 172094 333922 172162 333978
rect 172218 333922 202758 333978
rect 202814 333922 202882 333978
rect 202938 333922 233478 333978
rect 233534 333922 233602 333978
rect 233658 333922 264198 333978
rect 264254 333922 264322 333978
rect 264378 333922 285714 333978
rect 285770 333922 285838 333978
rect 285894 333922 285962 333978
rect 286018 333922 286086 333978
rect 286142 333922 301932 333978
rect 301988 333922 302056 333978
rect 302112 333922 302180 333978
rect 302236 333922 302304 333978
rect 302360 333922 316434 333978
rect 316490 333922 316558 333978
rect 316614 333922 316682 333978
rect 316738 333922 316806 333978
rect 316862 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 386614 333978
rect 386670 333922 386738 333978
rect 386794 333922 386862 333978
rect 386918 333922 386986 333978
rect 387042 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 499878 333978
rect 499934 333922 500002 333978
rect 500058 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect 277996 333658 475540 333674
rect 277996 333602 278012 333658
rect 278068 333602 475468 333658
rect 475524 333602 475540 333658
rect 277996 333586 475540 333602
rect 293228 332578 475540 332594
rect 293228 332522 293244 332578
rect 293300 332522 475468 332578
rect 475524 332522 475540 332578
rect 293228 332506 475540 332522
rect 299836 332398 475652 332414
rect 299836 332342 299852 332398
rect 299908 332342 475580 332398
rect 475636 332342 475652 332398
rect 299836 332326 475652 332342
rect 283036 330958 475540 330974
rect 283036 330902 283052 330958
rect 283108 330902 475468 330958
rect 475524 330902 475540 330958
rect 283036 330886 475540 330902
rect 273740 330058 352004 330074
rect 273740 330002 273756 330058
rect 273812 330002 351932 330058
rect 351988 330002 352004 330058
rect 273740 329986 352004 330002
rect 60156 329338 84996 329354
rect 60156 329282 60172 329338
rect 60228 329282 84924 329338
rect 84980 329282 84996 329338
rect 60156 329266 84996 329282
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 64518 328350
rect 64574 328294 64642 328350
rect 64698 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 95238 328350
rect 95294 328294 95362 328350
rect 95418 328294 125958 328350
rect 126014 328294 126082 328350
rect 126138 328294 156678 328350
rect 156734 328294 156802 328350
rect 156858 328294 187398 328350
rect 187454 328294 187522 328350
rect 187578 328294 218118 328350
rect 218174 328294 218242 328350
rect 218298 328294 248838 328350
rect 248894 328294 248962 328350
rect 249018 328294 281994 328350
rect 282050 328294 282118 328350
rect 282174 328294 282242 328350
rect 282298 328294 282366 328350
rect 282422 328294 302732 328350
rect 302788 328294 302856 328350
rect 302912 328294 302980 328350
rect 303036 328294 303104 328350
rect 303160 328294 312714 328350
rect 312770 328294 312838 328350
rect 312894 328294 312962 328350
rect 313018 328294 313086 328350
rect 313142 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 374154 328350
rect 374210 328294 374278 328350
rect 374334 328294 374402 328350
rect 374458 328294 374526 328350
rect 374582 328294 387414 328350
rect 387470 328294 387538 328350
rect 387594 328294 387662 328350
rect 387718 328294 387786 328350
rect 387842 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 484518 328350
rect 484574 328294 484642 328350
rect 484698 328294 515238 328350
rect 515294 328294 515362 328350
rect 515418 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 64518 328226
rect 64574 328170 64642 328226
rect 64698 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 95238 328226
rect 95294 328170 95362 328226
rect 95418 328170 125958 328226
rect 126014 328170 126082 328226
rect 126138 328170 156678 328226
rect 156734 328170 156802 328226
rect 156858 328170 187398 328226
rect 187454 328170 187522 328226
rect 187578 328170 218118 328226
rect 218174 328170 218242 328226
rect 218298 328170 248838 328226
rect 248894 328170 248962 328226
rect 249018 328170 281994 328226
rect 282050 328170 282118 328226
rect 282174 328170 282242 328226
rect 282298 328170 282366 328226
rect 282422 328170 302732 328226
rect 302788 328170 302856 328226
rect 302912 328170 302980 328226
rect 303036 328170 303104 328226
rect 303160 328170 312714 328226
rect 312770 328170 312838 328226
rect 312894 328170 312962 328226
rect 313018 328170 313086 328226
rect 313142 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 374154 328226
rect 374210 328170 374278 328226
rect 374334 328170 374402 328226
rect 374458 328170 374526 328226
rect 374582 328170 387414 328226
rect 387470 328170 387538 328226
rect 387594 328170 387662 328226
rect 387718 328170 387786 328226
rect 387842 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 484518 328226
rect 484574 328170 484642 328226
rect 484698 328170 515238 328226
rect 515294 328170 515362 328226
rect 515418 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 64518 328102
rect 64574 328046 64642 328102
rect 64698 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 95238 328102
rect 95294 328046 95362 328102
rect 95418 328046 125958 328102
rect 126014 328046 126082 328102
rect 126138 328046 156678 328102
rect 156734 328046 156802 328102
rect 156858 328046 187398 328102
rect 187454 328046 187522 328102
rect 187578 328046 218118 328102
rect 218174 328046 218242 328102
rect 218298 328046 248838 328102
rect 248894 328046 248962 328102
rect 249018 328046 281994 328102
rect 282050 328046 282118 328102
rect 282174 328046 282242 328102
rect 282298 328046 282366 328102
rect 282422 328046 302732 328102
rect 302788 328046 302856 328102
rect 302912 328046 302980 328102
rect 303036 328046 303104 328102
rect 303160 328046 312714 328102
rect 312770 328046 312838 328102
rect 312894 328046 312962 328102
rect 313018 328046 313086 328102
rect 313142 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 374154 328102
rect 374210 328046 374278 328102
rect 374334 328046 374402 328102
rect 374458 328046 374526 328102
rect 374582 328046 387414 328102
rect 387470 328046 387538 328102
rect 387594 328046 387662 328102
rect 387718 328046 387786 328102
rect 387842 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 484518 328102
rect 484574 328046 484642 328102
rect 484698 328046 515238 328102
rect 515294 328046 515362 328102
rect 515418 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 64518 327978
rect 64574 327922 64642 327978
rect 64698 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 95238 327978
rect 95294 327922 95362 327978
rect 95418 327922 125958 327978
rect 126014 327922 126082 327978
rect 126138 327922 156678 327978
rect 156734 327922 156802 327978
rect 156858 327922 187398 327978
rect 187454 327922 187522 327978
rect 187578 327922 218118 327978
rect 218174 327922 218242 327978
rect 218298 327922 248838 327978
rect 248894 327922 248962 327978
rect 249018 327922 281994 327978
rect 282050 327922 282118 327978
rect 282174 327922 282242 327978
rect 282298 327922 282366 327978
rect 282422 327922 302732 327978
rect 302788 327922 302856 327978
rect 302912 327922 302980 327978
rect 303036 327922 303104 327978
rect 303160 327922 312714 327978
rect 312770 327922 312838 327978
rect 312894 327922 312962 327978
rect 313018 327922 313086 327978
rect 313142 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 374154 327978
rect 374210 327922 374278 327978
rect 374334 327922 374402 327978
rect 374458 327922 374526 327978
rect 374582 327922 387414 327978
rect 387470 327922 387538 327978
rect 387594 327922 387662 327978
rect 387718 327922 387786 327978
rect 387842 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 484518 327978
rect 484574 327922 484642 327978
rect 484698 327922 515238 327978
rect 515294 327922 515362 327978
rect 515418 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect 60716 326818 74804 326834
rect 60716 326762 60732 326818
rect 60788 326762 74732 326818
rect 74788 326762 74804 326818
rect 60716 326746 74804 326762
rect 288300 326098 475540 326114
rect 288300 326042 288316 326098
rect 288372 326042 475468 326098
rect 475524 326042 475540 326098
rect 288300 326026 475540 326042
rect 273292 325018 353684 325034
rect 273292 324962 273308 325018
rect 273364 324962 353612 325018
rect 353668 324962 353684 325018
rect 273292 324946 353684 324962
rect 60380 324298 73124 324314
rect 60380 324242 60396 324298
rect 60452 324242 73052 324298
rect 73108 324242 73124 324298
rect 60380 324226 73124 324242
rect 273180 323398 360404 323414
rect 273180 323342 273196 323398
rect 273252 323342 360332 323398
rect 360388 323342 360404 323398
rect 273180 323326 360404 323342
rect 283036 321058 475540 321074
rect 283036 321002 283052 321058
rect 283108 321002 475468 321058
rect 475524 321002 475540 321058
rect 283036 320986 475540 321002
rect 272956 319978 348644 319994
rect 272956 319922 272972 319978
rect 273028 319922 348572 319978
rect 348628 319922 348644 319978
rect 272956 319906 348644 319922
rect 289868 317818 475540 317834
rect 289868 317762 289884 317818
rect 289940 317762 475468 317818
rect 475524 317762 475540 317818
rect 289868 317746 475540 317762
rect 274636 317638 475652 317654
rect 274636 317582 274652 317638
rect 274708 317582 475580 317638
rect 475636 317582 475652 317638
rect 274636 317566 475652 317582
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 79878 316350
rect 79934 316294 80002 316350
rect 80058 316294 110598 316350
rect 110654 316294 110722 316350
rect 110778 316294 141318 316350
rect 141374 316294 141442 316350
rect 141498 316294 172038 316350
rect 172094 316294 172162 316350
rect 172218 316294 202758 316350
rect 202814 316294 202882 316350
rect 202938 316294 233478 316350
rect 233534 316294 233602 316350
rect 233658 316294 264198 316350
rect 264254 316294 264322 316350
rect 264378 316294 285714 316350
rect 285770 316294 285838 316350
rect 285894 316294 285962 316350
rect 286018 316294 286086 316350
rect 286142 316294 301932 316350
rect 301988 316294 302056 316350
rect 302112 316294 302180 316350
rect 302236 316294 302304 316350
rect 302360 316294 316434 316350
rect 316490 316294 316558 316350
rect 316614 316294 316682 316350
rect 316738 316294 316806 316350
rect 316862 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 386614 316350
rect 386670 316294 386738 316350
rect 386794 316294 386862 316350
rect 386918 316294 386986 316350
rect 387042 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 499878 316350
rect 499934 316294 500002 316350
rect 500058 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 79878 316226
rect 79934 316170 80002 316226
rect 80058 316170 110598 316226
rect 110654 316170 110722 316226
rect 110778 316170 141318 316226
rect 141374 316170 141442 316226
rect 141498 316170 172038 316226
rect 172094 316170 172162 316226
rect 172218 316170 202758 316226
rect 202814 316170 202882 316226
rect 202938 316170 233478 316226
rect 233534 316170 233602 316226
rect 233658 316170 264198 316226
rect 264254 316170 264322 316226
rect 264378 316170 285714 316226
rect 285770 316170 285838 316226
rect 285894 316170 285962 316226
rect 286018 316170 286086 316226
rect 286142 316170 301932 316226
rect 301988 316170 302056 316226
rect 302112 316170 302180 316226
rect 302236 316170 302304 316226
rect 302360 316170 316434 316226
rect 316490 316170 316558 316226
rect 316614 316170 316682 316226
rect 316738 316170 316806 316226
rect 316862 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 386614 316226
rect 386670 316170 386738 316226
rect 386794 316170 386862 316226
rect 386918 316170 386986 316226
rect 387042 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 499878 316226
rect 499934 316170 500002 316226
rect 500058 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 79878 316102
rect 79934 316046 80002 316102
rect 80058 316046 110598 316102
rect 110654 316046 110722 316102
rect 110778 316046 141318 316102
rect 141374 316046 141442 316102
rect 141498 316046 172038 316102
rect 172094 316046 172162 316102
rect 172218 316046 202758 316102
rect 202814 316046 202882 316102
rect 202938 316046 233478 316102
rect 233534 316046 233602 316102
rect 233658 316046 264198 316102
rect 264254 316046 264322 316102
rect 264378 316046 285714 316102
rect 285770 316046 285838 316102
rect 285894 316046 285962 316102
rect 286018 316046 286086 316102
rect 286142 316046 301932 316102
rect 301988 316046 302056 316102
rect 302112 316046 302180 316102
rect 302236 316046 302304 316102
rect 302360 316046 316434 316102
rect 316490 316046 316558 316102
rect 316614 316046 316682 316102
rect 316738 316046 316806 316102
rect 316862 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 386614 316102
rect 386670 316046 386738 316102
rect 386794 316046 386862 316102
rect 386918 316046 386986 316102
rect 387042 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 499878 316102
rect 499934 316046 500002 316102
rect 500058 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 79878 315978
rect 79934 315922 80002 315978
rect 80058 315922 110598 315978
rect 110654 315922 110722 315978
rect 110778 315922 141318 315978
rect 141374 315922 141442 315978
rect 141498 315922 172038 315978
rect 172094 315922 172162 315978
rect 172218 315922 202758 315978
rect 202814 315922 202882 315978
rect 202938 315922 233478 315978
rect 233534 315922 233602 315978
rect 233658 315922 264198 315978
rect 264254 315922 264322 315978
rect 264378 315922 285714 315978
rect 285770 315922 285838 315978
rect 285894 315922 285962 315978
rect 286018 315922 286086 315978
rect 286142 315922 301932 315978
rect 301988 315922 302056 315978
rect 302112 315922 302180 315978
rect 302236 315922 302304 315978
rect 302360 315922 316434 315978
rect 316490 315922 316558 315978
rect 316614 315922 316682 315978
rect 316738 315922 316806 315978
rect 316862 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 386614 315978
rect 386670 315922 386738 315978
rect 386794 315922 386862 315978
rect 386918 315922 386986 315978
rect 387042 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 499878 315978
rect 499934 315922 500002 315978
rect 500058 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect 293228 314218 475540 314234
rect 293228 314162 293244 314218
rect 293300 314162 475468 314218
rect 475524 314162 475540 314218
rect 293228 314146 475540 314162
rect 281356 312598 475540 312614
rect 281356 312542 281372 312598
rect 281428 312542 475468 312598
rect 475524 312542 475540 312598
rect 281356 312526 475540 312542
rect 273068 311698 350324 311714
rect 273068 311642 273084 311698
rect 273140 311642 350252 311698
rect 350308 311642 350324 311698
rect 273068 311626 350324 311642
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 64518 310350
rect 64574 310294 64642 310350
rect 64698 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 95238 310350
rect 95294 310294 95362 310350
rect 95418 310294 125958 310350
rect 126014 310294 126082 310350
rect 126138 310294 156678 310350
rect 156734 310294 156802 310350
rect 156858 310294 187398 310350
rect 187454 310294 187522 310350
rect 187578 310294 218118 310350
rect 218174 310294 218242 310350
rect 218298 310294 248838 310350
rect 248894 310294 248962 310350
rect 249018 310294 281994 310350
rect 282050 310294 282118 310350
rect 282174 310294 282242 310350
rect 282298 310294 282366 310350
rect 282422 310294 302732 310350
rect 302788 310294 302856 310350
rect 302912 310294 302980 310350
rect 303036 310294 303104 310350
rect 303160 310294 312714 310350
rect 312770 310294 312838 310350
rect 312894 310294 312962 310350
rect 313018 310294 313086 310350
rect 313142 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 374154 310350
rect 374210 310294 374278 310350
rect 374334 310294 374402 310350
rect 374458 310294 374526 310350
rect 374582 310294 387414 310350
rect 387470 310294 387538 310350
rect 387594 310294 387662 310350
rect 387718 310294 387786 310350
rect 387842 310294 404874 310350
rect 404930 310294 404998 310350
rect 405054 310294 405122 310350
rect 405178 310294 405246 310350
rect 405302 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 484518 310350
rect 484574 310294 484642 310350
rect 484698 310294 515238 310350
rect 515294 310294 515362 310350
rect 515418 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 64518 310226
rect 64574 310170 64642 310226
rect 64698 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 95238 310226
rect 95294 310170 95362 310226
rect 95418 310170 125958 310226
rect 126014 310170 126082 310226
rect 126138 310170 156678 310226
rect 156734 310170 156802 310226
rect 156858 310170 187398 310226
rect 187454 310170 187522 310226
rect 187578 310170 218118 310226
rect 218174 310170 218242 310226
rect 218298 310170 248838 310226
rect 248894 310170 248962 310226
rect 249018 310170 281994 310226
rect 282050 310170 282118 310226
rect 282174 310170 282242 310226
rect 282298 310170 282366 310226
rect 282422 310170 302732 310226
rect 302788 310170 302856 310226
rect 302912 310170 302980 310226
rect 303036 310170 303104 310226
rect 303160 310170 312714 310226
rect 312770 310170 312838 310226
rect 312894 310170 312962 310226
rect 313018 310170 313086 310226
rect 313142 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 374154 310226
rect 374210 310170 374278 310226
rect 374334 310170 374402 310226
rect 374458 310170 374526 310226
rect 374582 310170 387414 310226
rect 387470 310170 387538 310226
rect 387594 310170 387662 310226
rect 387718 310170 387786 310226
rect 387842 310170 404874 310226
rect 404930 310170 404998 310226
rect 405054 310170 405122 310226
rect 405178 310170 405246 310226
rect 405302 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 484518 310226
rect 484574 310170 484642 310226
rect 484698 310170 515238 310226
rect 515294 310170 515362 310226
rect 515418 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 64518 310102
rect 64574 310046 64642 310102
rect 64698 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 95238 310102
rect 95294 310046 95362 310102
rect 95418 310046 125958 310102
rect 126014 310046 126082 310102
rect 126138 310046 156678 310102
rect 156734 310046 156802 310102
rect 156858 310046 187398 310102
rect 187454 310046 187522 310102
rect 187578 310046 218118 310102
rect 218174 310046 218242 310102
rect 218298 310046 248838 310102
rect 248894 310046 248962 310102
rect 249018 310046 281994 310102
rect 282050 310046 282118 310102
rect 282174 310046 282242 310102
rect 282298 310046 282366 310102
rect 282422 310046 302732 310102
rect 302788 310046 302856 310102
rect 302912 310046 302980 310102
rect 303036 310046 303104 310102
rect 303160 310046 312714 310102
rect 312770 310046 312838 310102
rect 312894 310046 312962 310102
rect 313018 310046 313086 310102
rect 313142 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 374154 310102
rect 374210 310046 374278 310102
rect 374334 310046 374402 310102
rect 374458 310046 374526 310102
rect 374582 310046 387414 310102
rect 387470 310046 387538 310102
rect 387594 310046 387662 310102
rect 387718 310046 387786 310102
rect 387842 310046 404874 310102
rect 404930 310046 404998 310102
rect 405054 310046 405122 310102
rect 405178 310046 405246 310102
rect 405302 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 484518 310102
rect 484574 310046 484642 310102
rect 484698 310046 515238 310102
rect 515294 310046 515362 310102
rect 515418 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 64518 309978
rect 64574 309922 64642 309978
rect 64698 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 95238 309978
rect 95294 309922 95362 309978
rect 95418 309922 125958 309978
rect 126014 309922 126082 309978
rect 126138 309922 156678 309978
rect 156734 309922 156802 309978
rect 156858 309922 187398 309978
rect 187454 309922 187522 309978
rect 187578 309922 218118 309978
rect 218174 309922 218242 309978
rect 218298 309922 248838 309978
rect 248894 309922 248962 309978
rect 249018 309922 281994 309978
rect 282050 309922 282118 309978
rect 282174 309922 282242 309978
rect 282298 309922 282366 309978
rect 282422 309922 302732 309978
rect 302788 309922 302856 309978
rect 302912 309922 302980 309978
rect 303036 309922 303104 309978
rect 303160 309922 312714 309978
rect 312770 309922 312838 309978
rect 312894 309922 312962 309978
rect 313018 309922 313086 309978
rect 313142 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 374154 309978
rect 374210 309922 374278 309978
rect 374334 309922 374402 309978
rect 374458 309922 374526 309978
rect 374582 309922 387414 309978
rect 387470 309922 387538 309978
rect 387594 309922 387662 309978
rect 387718 309922 387786 309978
rect 387842 309922 404874 309978
rect 404930 309922 404998 309978
rect 405054 309922 405122 309978
rect 405178 309922 405246 309978
rect 405302 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 484518 309978
rect 484574 309922 484642 309978
rect 484698 309922 515238 309978
rect 515294 309922 515362 309978
rect 515418 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect 60716 307558 76596 307574
rect 60716 307502 60732 307558
rect 60788 307502 76524 307558
rect 76580 307502 76596 307558
rect 60716 307486 76596 307502
rect 276316 307558 475540 307574
rect 276316 307502 276332 307558
rect 276388 307502 475468 307558
rect 475524 307502 475540 307558
rect 276316 307486 475540 307502
rect 57916 301798 388068 301814
rect 57916 301742 57932 301798
rect 57988 301742 387996 301798
rect 388052 301742 388068 301798
rect 57916 301726 388068 301742
rect 60492 301618 590900 301634
rect 60492 301562 60508 301618
rect 60564 301562 590828 301618
rect 590884 301562 590900 301618
rect 60492 301546 590900 301562
rect 53100 300718 591012 300734
rect 53100 300662 53116 300718
rect 53172 300662 590940 300718
rect 590996 300662 591012 300718
rect 53100 300646 591012 300662
rect 4156 300538 474644 300554
rect 4156 300482 4172 300538
rect 4228 300482 474572 300538
rect 474628 300482 474644 300538
rect 4156 300466 474644 300482
rect 54332 300358 388068 300374
rect 54332 300302 54348 300358
rect 54404 300302 387996 300358
rect 388052 300302 388068 300358
rect 54332 300286 388068 300302
rect 388204 300358 388292 300374
rect 388204 300302 388220 300358
rect 388276 300302 388292 300358
rect 388204 300194 388292 300302
rect 84796 300178 388292 300194
rect 84796 300122 84812 300178
rect 84868 300122 388292 300178
rect 84796 300106 388292 300122
rect 83788 298918 480244 298934
rect 83788 298862 83804 298918
rect 83860 298862 480172 298918
rect 480228 298862 480244 298918
rect 83788 298846 480244 298862
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 79878 298350
rect 79934 298294 80002 298350
rect 80058 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 110598 298350
rect 110654 298294 110722 298350
rect 110778 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 141318 298350
rect 141374 298294 141442 298350
rect 141498 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 172038 298350
rect 172094 298294 172162 298350
rect 172218 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 202758 298350
rect 202814 298294 202882 298350
rect 202938 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 233478 298350
rect 233534 298294 233602 298350
rect 233658 298294 254994 298350
rect 255050 298294 255118 298350
rect 255174 298294 255242 298350
rect 255298 298294 255366 298350
rect 255422 298294 264198 298350
rect 264254 298294 264322 298350
rect 264378 298294 285714 298350
rect 285770 298294 285838 298350
rect 285894 298294 285962 298350
rect 286018 298294 286086 298350
rect 286142 298294 301932 298350
rect 301988 298294 302056 298350
rect 302112 298294 302180 298350
rect 302236 298294 302304 298350
rect 302360 298294 316434 298350
rect 316490 298294 316558 298350
rect 316614 298294 316682 298350
rect 316738 298294 316806 298350
rect 316862 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 386614 298350
rect 386670 298294 386738 298350
rect 386794 298294 386862 298350
rect 386918 298294 386986 298350
rect 387042 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 79878 298226
rect 79934 298170 80002 298226
rect 80058 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 110598 298226
rect 110654 298170 110722 298226
rect 110778 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 141318 298226
rect 141374 298170 141442 298226
rect 141498 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 172038 298226
rect 172094 298170 172162 298226
rect 172218 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 202758 298226
rect 202814 298170 202882 298226
rect 202938 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 233478 298226
rect 233534 298170 233602 298226
rect 233658 298170 254994 298226
rect 255050 298170 255118 298226
rect 255174 298170 255242 298226
rect 255298 298170 255366 298226
rect 255422 298170 264198 298226
rect 264254 298170 264322 298226
rect 264378 298170 285714 298226
rect 285770 298170 285838 298226
rect 285894 298170 285962 298226
rect 286018 298170 286086 298226
rect 286142 298170 301932 298226
rect 301988 298170 302056 298226
rect 302112 298170 302180 298226
rect 302236 298170 302304 298226
rect 302360 298170 316434 298226
rect 316490 298170 316558 298226
rect 316614 298170 316682 298226
rect 316738 298170 316806 298226
rect 316862 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 386614 298226
rect 386670 298170 386738 298226
rect 386794 298170 386862 298226
rect 386918 298170 386986 298226
rect 387042 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 79878 298102
rect 79934 298046 80002 298102
rect 80058 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 110598 298102
rect 110654 298046 110722 298102
rect 110778 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 141318 298102
rect 141374 298046 141442 298102
rect 141498 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 172038 298102
rect 172094 298046 172162 298102
rect 172218 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 202758 298102
rect 202814 298046 202882 298102
rect 202938 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 233478 298102
rect 233534 298046 233602 298102
rect 233658 298046 254994 298102
rect 255050 298046 255118 298102
rect 255174 298046 255242 298102
rect 255298 298046 255366 298102
rect 255422 298046 264198 298102
rect 264254 298046 264322 298102
rect 264378 298046 285714 298102
rect 285770 298046 285838 298102
rect 285894 298046 285962 298102
rect 286018 298046 286086 298102
rect 286142 298046 301932 298102
rect 301988 298046 302056 298102
rect 302112 298046 302180 298102
rect 302236 298046 302304 298102
rect 302360 298046 316434 298102
rect 316490 298046 316558 298102
rect 316614 298046 316682 298102
rect 316738 298046 316806 298102
rect 316862 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 386614 298102
rect 386670 298046 386738 298102
rect 386794 298046 386862 298102
rect 386918 298046 386986 298102
rect 387042 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 79878 297978
rect 79934 297922 80002 297978
rect 80058 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 110598 297978
rect 110654 297922 110722 297978
rect 110778 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 141318 297978
rect 141374 297922 141442 297978
rect 141498 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 172038 297978
rect 172094 297922 172162 297978
rect 172218 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 202758 297978
rect 202814 297922 202882 297978
rect 202938 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 233478 297978
rect 233534 297922 233602 297978
rect 233658 297922 254994 297978
rect 255050 297922 255118 297978
rect 255174 297922 255242 297978
rect 255298 297922 255366 297978
rect 255422 297922 264198 297978
rect 264254 297922 264322 297978
rect 264378 297922 285714 297978
rect 285770 297922 285838 297978
rect 285894 297922 285962 297978
rect 286018 297922 286086 297978
rect 286142 297922 301932 297978
rect 301988 297922 302056 297978
rect 302112 297922 302180 297978
rect 302236 297922 302304 297978
rect 302360 297922 316434 297978
rect 316490 297922 316558 297978
rect 316614 297922 316682 297978
rect 316738 297922 316806 297978
rect 316862 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 386614 297978
rect 386670 297922 386738 297978
rect 386794 297922 386862 297978
rect 386918 297922 386986 297978
rect 387042 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect 84908 297298 591124 297314
rect 84908 297242 84924 297298
rect 84980 297242 591052 297298
rect 591108 297242 591124 297298
rect 84908 297226 591124 297242
rect 56908 297118 390644 297134
rect 56908 297062 56924 297118
rect 56980 297062 390572 297118
rect 390628 297062 390644 297118
rect 56908 297046 390644 297062
rect 53548 296938 388516 296954
rect 53548 296882 53564 296938
rect 53620 296882 388444 296938
rect 388500 296882 388516 296938
rect 53548 296866 388516 296882
rect 58476 296758 388068 296774
rect 58476 296702 58492 296758
rect 58548 296702 387996 296758
rect 388052 296702 388068 296758
rect 58476 296686 388068 296702
rect 58140 295678 591348 295694
rect 58140 295622 58156 295678
rect 58212 295622 591276 295678
rect 591332 295622 591348 295678
rect 58140 295606 591348 295622
rect 58700 295498 590564 295514
rect 58700 295442 58716 295498
rect 58772 295442 590492 295498
rect 590548 295442 590564 295498
rect 58700 295426 590564 295442
rect 83564 295318 480020 295334
rect 83564 295262 83580 295318
rect 83636 295262 479948 295318
rect 480004 295262 480020 295318
rect 83564 295246 480020 295262
rect 83676 295138 479796 295154
rect 83676 295082 83692 295138
rect 83748 295082 479724 295138
rect 479780 295082 479796 295138
rect 83676 295066 479796 295082
rect 4268 293878 480132 293894
rect 4268 293822 4284 293878
rect 4340 293822 480060 293878
rect 480116 293822 480132 293878
rect 4268 293806 480132 293822
rect 53212 293698 476996 293714
rect 53212 293642 53228 293698
rect 53284 293642 476924 293698
rect 476980 293642 476996 293698
rect 53212 293626 476996 293642
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 251274 292350
rect 251330 292294 251398 292350
rect 251454 292294 251522 292350
rect 251578 292294 251646 292350
rect 251702 292294 281994 292350
rect 282050 292294 282118 292350
rect 282174 292294 282242 292350
rect 282298 292294 282366 292350
rect 282422 292294 302732 292350
rect 302788 292294 302856 292350
rect 302912 292294 302980 292350
rect 303036 292294 303104 292350
rect 303160 292294 312714 292350
rect 312770 292294 312838 292350
rect 312894 292294 312962 292350
rect 313018 292294 313086 292350
rect 313142 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 374154 292350
rect 374210 292294 374278 292350
rect 374334 292294 374402 292350
rect 374458 292294 374526 292350
rect 374582 292294 387414 292350
rect 387470 292294 387538 292350
rect 387594 292294 387662 292350
rect 387718 292294 387786 292350
rect 387842 292294 404874 292350
rect 404930 292294 404998 292350
rect 405054 292294 405122 292350
rect 405178 292294 405246 292350
rect 405302 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 251274 292226
rect 251330 292170 251398 292226
rect 251454 292170 251522 292226
rect 251578 292170 251646 292226
rect 251702 292170 281994 292226
rect 282050 292170 282118 292226
rect 282174 292170 282242 292226
rect 282298 292170 282366 292226
rect 282422 292170 302732 292226
rect 302788 292170 302856 292226
rect 302912 292170 302980 292226
rect 303036 292170 303104 292226
rect 303160 292170 312714 292226
rect 312770 292170 312838 292226
rect 312894 292170 312962 292226
rect 313018 292170 313086 292226
rect 313142 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 374154 292226
rect 374210 292170 374278 292226
rect 374334 292170 374402 292226
rect 374458 292170 374526 292226
rect 374582 292170 387414 292226
rect 387470 292170 387538 292226
rect 387594 292170 387662 292226
rect 387718 292170 387786 292226
rect 387842 292170 404874 292226
rect 404930 292170 404998 292226
rect 405054 292170 405122 292226
rect 405178 292170 405246 292226
rect 405302 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 251274 292102
rect 251330 292046 251398 292102
rect 251454 292046 251522 292102
rect 251578 292046 251646 292102
rect 251702 292046 281994 292102
rect 282050 292046 282118 292102
rect 282174 292046 282242 292102
rect 282298 292046 282366 292102
rect 282422 292046 302732 292102
rect 302788 292046 302856 292102
rect 302912 292046 302980 292102
rect 303036 292046 303104 292102
rect 303160 292046 312714 292102
rect 312770 292046 312838 292102
rect 312894 292046 312962 292102
rect 313018 292046 313086 292102
rect 313142 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 374154 292102
rect 374210 292046 374278 292102
rect 374334 292046 374402 292102
rect 374458 292046 374526 292102
rect 374582 292046 387414 292102
rect 387470 292046 387538 292102
rect 387594 292046 387662 292102
rect 387718 292046 387786 292102
rect 387842 292046 404874 292102
rect 404930 292046 404998 292102
rect 405054 292046 405122 292102
rect 405178 292046 405246 292102
rect 405302 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 251274 291978
rect 251330 291922 251398 291978
rect 251454 291922 251522 291978
rect 251578 291922 251646 291978
rect 251702 291922 281994 291978
rect 282050 291922 282118 291978
rect 282174 291922 282242 291978
rect 282298 291922 282366 291978
rect 282422 291922 302732 291978
rect 302788 291922 302856 291978
rect 302912 291922 302980 291978
rect 303036 291922 303104 291978
rect 303160 291922 312714 291978
rect 312770 291922 312838 291978
rect 312894 291922 312962 291978
rect 313018 291922 313086 291978
rect 313142 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 374154 291978
rect 374210 291922 374278 291978
rect 374334 291922 374402 291978
rect 374458 291922 374526 291978
rect 374582 291922 387414 291978
rect 387470 291922 387538 291978
rect 387594 291922 387662 291978
rect 387718 291922 387786 291978
rect 387842 291922 404874 291978
rect 404930 291922 404998 291978
rect 405054 291922 405122 291978
rect 405178 291922 405246 291978
rect 405302 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect 53660 291718 388068 291734
rect 53660 291662 53676 291718
rect 53732 291662 387996 291718
rect 388052 291662 388068 291718
rect 53660 291646 388068 291662
rect 54780 290638 476212 290654
rect 54780 290582 54796 290638
rect 54852 290582 476140 290638
rect 476196 290582 476212 290638
rect 54780 290566 476212 290582
rect 69676 290458 476772 290474
rect 69676 290402 69692 290458
rect 69748 290402 476700 290458
rect 476756 290402 476772 290458
rect 69676 290386 476772 290402
rect 55004 290278 388068 290294
rect 55004 290222 55020 290278
rect 55076 290222 387996 290278
rect 388052 290222 388068 290278
rect 55004 290206 388068 290222
rect 60268 288838 591236 288854
rect 60268 288782 60284 288838
rect 60340 288782 591164 288838
rect 591220 288782 591236 288838
rect 60268 288766 591236 288782
rect 4380 288658 478228 288674
rect 4380 288602 4396 288658
rect 4452 288602 478156 288658
rect 478212 288602 478228 288658
rect 4380 288586 478228 288602
rect 54556 288478 476100 288494
rect 54556 288422 54572 288478
rect 54628 288422 476028 288478
rect 476084 288422 476100 288478
rect 54556 288406 476100 288422
rect 53436 287218 476660 287234
rect 53436 287162 53452 287218
rect 53508 287162 476588 287218
rect 476644 287162 476660 287218
rect 53436 287146 476660 287162
rect 60156 287038 476884 287054
rect 60156 286982 60172 287038
rect 60228 286982 476812 287038
rect 476868 286982 476884 287038
rect 60156 286966 476884 286982
rect 78076 286858 477108 286874
rect 78076 286802 78092 286858
rect 78148 286802 477036 286858
rect 477092 286802 477108 286858
rect 78076 286786 477108 286802
rect 76508 285598 590788 285614
rect 76508 285542 76524 285598
rect 76580 285542 590716 285598
rect 590772 285542 590788 285598
rect 76508 285526 590788 285542
rect 53324 285418 476436 285434
rect 53324 285362 53340 285418
rect 53396 285362 476364 285418
rect 476420 285362 476436 285418
rect 53324 285346 476436 285362
rect 291548 285238 590228 285254
rect 291548 285182 291564 285238
rect 291620 285182 590156 285238
rect 590212 285182 590228 285238
rect 291548 285166 590228 285182
rect 4940 283798 479908 283814
rect 4940 283742 4956 283798
rect 5012 283742 479836 283798
rect 479892 283742 479908 283798
rect 4940 283726 479908 283742
rect 60044 283618 475540 283634
rect 60044 283562 60060 283618
rect 60116 283562 475468 283618
rect 475524 283562 475540 283618
rect 60044 283546 475540 283562
rect 55116 282178 590900 282194
rect 55116 282122 55132 282178
rect 55188 282122 590828 282178
rect 590884 282122 590900 282178
rect 55116 282106 590900 282122
rect 58588 281998 590676 282014
rect 58588 281942 58604 281998
rect 58660 281942 590604 281998
rect 590660 281942 590676 281998
rect 58588 281926 590676 281942
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 70674 280350
rect 70730 280294 70798 280350
rect 70854 280294 70922 280350
rect 70978 280294 71046 280350
rect 71102 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 254994 280350
rect 255050 280294 255118 280350
rect 255174 280294 255242 280350
rect 255298 280294 255366 280350
rect 255422 280294 285714 280350
rect 285770 280294 285838 280350
rect 285894 280294 285962 280350
rect 286018 280294 286086 280350
rect 286142 280294 316434 280350
rect 316490 280294 316558 280350
rect 316614 280294 316682 280350
rect 316738 280294 316806 280350
rect 316862 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 408594 280350
rect 408650 280294 408718 280350
rect 408774 280294 408842 280350
rect 408898 280294 408966 280350
rect 409022 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 70674 280226
rect 70730 280170 70798 280226
rect 70854 280170 70922 280226
rect 70978 280170 71046 280226
rect 71102 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 254994 280226
rect 255050 280170 255118 280226
rect 255174 280170 255242 280226
rect 255298 280170 255366 280226
rect 255422 280170 285714 280226
rect 285770 280170 285838 280226
rect 285894 280170 285962 280226
rect 286018 280170 286086 280226
rect 286142 280170 316434 280226
rect 316490 280170 316558 280226
rect 316614 280170 316682 280226
rect 316738 280170 316806 280226
rect 316862 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 408594 280226
rect 408650 280170 408718 280226
rect 408774 280170 408842 280226
rect 408898 280170 408966 280226
rect 409022 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 70674 280102
rect 70730 280046 70798 280102
rect 70854 280046 70922 280102
rect 70978 280046 71046 280102
rect 71102 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 254994 280102
rect 255050 280046 255118 280102
rect 255174 280046 255242 280102
rect 255298 280046 255366 280102
rect 255422 280046 285714 280102
rect 285770 280046 285838 280102
rect 285894 280046 285962 280102
rect 286018 280046 286086 280102
rect 286142 280046 316434 280102
rect 316490 280046 316558 280102
rect 316614 280046 316682 280102
rect 316738 280046 316806 280102
rect 316862 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 408594 280102
rect 408650 280046 408718 280102
rect 408774 280046 408842 280102
rect 408898 280046 408966 280102
rect 409022 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 70674 279978
rect 70730 279922 70798 279978
rect 70854 279922 70922 279978
rect 70978 279922 71046 279978
rect 71102 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 254994 279978
rect 255050 279922 255118 279978
rect 255174 279922 255242 279978
rect 255298 279922 255366 279978
rect 255422 279922 285714 279978
rect 285770 279922 285838 279978
rect 285894 279922 285962 279978
rect 286018 279922 286086 279978
rect 286142 279922 316434 279978
rect 316490 279922 316558 279978
rect 316614 279922 316682 279978
rect 316738 279922 316806 279978
rect 316862 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 408594 279978
rect 408650 279922 408718 279978
rect 408774 279922 408842 279978
rect 408898 279922 408966 279978
rect 409022 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 66954 274350
rect 67010 274294 67078 274350
rect 67134 274294 67202 274350
rect 67258 274294 67326 274350
rect 67382 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 251274 274350
rect 251330 274294 251398 274350
rect 251454 274294 251522 274350
rect 251578 274294 251646 274350
rect 251702 274294 281994 274350
rect 282050 274294 282118 274350
rect 282174 274294 282242 274350
rect 282298 274294 282366 274350
rect 282422 274294 312714 274350
rect 312770 274294 312838 274350
rect 312894 274294 312962 274350
rect 313018 274294 313086 274350
rect 313142 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 374154 274350
rect 374210 274294 374278 274350
rect 374334 274294 374402 274350
rect 374458 274294 374526 274350
rect 374582 274294 404874 274350
rect 404930 274294 404998 274350
rect 405054 274294 405122 274350
rect 405178 274294 405246 274350
rect 405302 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 66954 274226
rect 67010 274170 67078 274226
rect 67134 274170 67202 274226
rect 67258 274170 67326 274226
rect 67382 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 251274 274226
rect 251330 274170 251398 274226
rect 251454 274170 251522 274226
rect 251578 274170 251646 274226
rect 251702 274170 281994 274226
rect 282050 274170 282118 274226
rect 282174 274170 282242 274226
rect 282298 274170 282366 274226
rect 282422 274170 312714 274226
rect 312770 274170 312838 274226
rect 312894 274170 312962 274226
rect 313018 274170 313086 274226
rect 313142 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 374154 274226
rect 374210 274170 374278 274226
rect 374334 274170 374402 274226
rect 374458 274170 374526 274226
rect 374582 274170 404874 274226
rect 404930 274170 404998 274226
rect 405054 274170 405122 274226
rect 405178 274170 405246 274226
rect 405302 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 66954 274102
rect 67010 274046 67078 274102
rect 67134 274046 67202 274102
rect 67258 274046 67326 274102
rect 67382 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 251274 274102
rect 251330 274046 251398 274102
rect 251454 274046 251522 274102
rect 251578 274046 251646 274102
rect 251702 274046 281994 274102
rect 282050 274046 282118 274102
rect 282174 274046 282242 274102
rect 282298 274046 282366 274102
rect 282422 274046 312714 274102
rect 312770 274046 312838 274102
rect 312894 274046 312962 274102
rect 313018 274046 313086 274102
rect 313142 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 374154 274102
rect 374210 274046 374278 274102
rect 374334 274046 374402 274102
rect 374458 274046 374526 274102
rect 374582 274046 404874 274102
rect 404930 274046 404998 274102
rect 405054 274046 405122 274102
rect 405178 274046 405246 274102
rect 405302 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 66954 273978
rect 67010 273922 67078 273978
rect 67134 273922 67202 273978
rect 67258 273922 67326 273978
rect 67382 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 251274 273978
rect 251330 273922 251398 273978
rect 251454 273922 251522 273978
rect 251578 273922 251646 273978
rect 251702 273922 281994 273978
rect 282050 273922 282118 273978
rect 282174 273922 282242 273978
rect 282298 273922 282366 273978
rect 282422 273922 312714 273978
rect 312770 273922 312838 273978
rect 312894 273922 312962 273978
rect 313018 273922 313086 273978
rect 313142 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 374154 273978
rect 374210 273922 374278 273978
rect 374334 273922 374402 273978
rect 374458 273922 374526 273978
rect 374582 273922 404874 273978
rect 404930 273922 404998 273978
rect 405054 273922 405122 273978
rect 405178 273922 405246 273978
rect 405302 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 70674 262350
rect 70730 262294 70798 262350
rect 70854 262294 70922 262350
rect 70978 262294 71046 262350
rect 71102 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 254994 262350
rect 255050 262294 255118 262350
rect 255174 262294 255242 262350
rect 255298 262294 255366 262350
rect 255422 262294 285714 262350
rect 285770 262294 285838 262350
rect 285894 262294 285962 262350
rect 286018 262294 286086 262350
rect 286142 262294 316434 262350
rect 316490 262294 316558 262350
rect 316614 262294 316682 262350
rect 316738 262294 316806 262350
rect 316862 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 70674 262226
rect 70730 262170 70798 262226
rect 70854 262170 70922 262226
rect 70978 262170 71046 262226
rect 71102 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 254994 262226
rect 255050 262170 255118 262226
rect 255174 262170 255242 262226
rect 255298 262170 255366 262226
rect 255422 262170 285714 262226
rect 285770 262170 285838 262226
rect 285894 262170 285962 262226
rect 286018 262170 286086 262226
rect 286142 262170 316434 262226
rect 316490 262170 316558 262226
rect 316614 262170 316682 262226
rect 316738 262170 316806 262226
rect 316862 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 70674 262102
rect 70730 262046 70798 262102
rect 70854 262046 70922 262102
rect 70978 262046 71046 262102
rect 71102 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 254994 262102
rect 255050 262046 255118 262102
rect 255174 262046 255242 262102
rect 255298 262046 255366 262102
rect 255422 262046 285714 262102
rect 285770 262046 285838 262102
rect 285894 262046 285962 262102
rect 286018 262046 286086 262102
rect 286142 262046 316434 262102
rect 316490 262046 316558 262102
rect 316614 262046 316682 262102
rect 316738 262046 316806 262102
rect 316862 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 70674 261978
rect 70730 261922 70798 261978
rect 70854 261922 70922 261978
rect 70978 261922 71046 261978
rect 71102 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 254994 261978
rect 255050 261922 255118 261978
rect 255174 261922 255242 261978
rect 255298 261922 255366 261978
rect 255422 261922 285714 261978
rect 285770 261922 285838 261978
rect 285894 261922 285962 261978
rect 286018 261922 286086 261978
rect 286142 261922 316434 261978
rect 316490 261922 316558 261978
rect 316614 261922 316682 261978
rect 316738 261922 316806 261978
rect 316862 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 66954 256350
rect 67010 256294 67078 256350
rect 67134 256294 67202 256350
rect 67258 256294 67326 256350
rect 67382 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 251274 256350
rect 251330 256294 251398 256350
rect 251454 256294 251522 256350
rect 251578 256294 251646 256350
rect 251702 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 404874 256350
rect 404930 256294 404998 256350
rect 405054 256294 405122 256350
rect 405178 256294 405246 256350
rect 405302 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 66954 256226
rect 67010 256170 67078 256226
rect 67134 256170 67202 256226
rect 67258 256170 67326 256226
rect 67382 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 251274 256226
rect 251330 256170 251398 256226
rect 251454 256170 251522 256226
rect 251578 256170 251646 256226
rect 251702 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 404874 256226
rect 404930 256170 404998 256226
rect 405054 256170 405122 256226
rect 405178 256170 405246 256226
rect 405302 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 66954 256102
rect 67010 256046 67078 256102
rect 67134 256046 67202 256102
rect 67258 256046 67326 256102
rect 67382 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 251274 256102
rect 251330 256046 251398 256102
rect 251454 256046 251522 256102
rect 251578 256046 251646 256102
rect 251702 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 404874 256102
rect 404930 256046 404998 256102
rect 405054 256046 405122 256102
rect 405178 256046 405246 256102
rect 405302 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 256023 597980 256046
rect -1916 255978 472732 256023
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 66954 255978
rect 67010 255922 67078 255978
rect 67134 255922 67202 255978
rect 67258 255922 67326 255978
rect 67382 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 251274 255978
rect 251330 255922 251398 255978
rect 251454 255922 251522 255978
rect 251578 255922 251646 255978
rect 251702 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 404874 255978
rect 404930 255922 404998 255978
rect 405054 255922 405122 255978
rect 405178 255922 405246 255978
rect 405302 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255967 472732 255978
rect 472788 255967 472856 256023
rect 472912 255967 472980 256023
rect 473036 255967 473104 256023
rect 473160 255978 557414 256023
rect 473160 255967 497034 255978
rect 466742 255922 497034 255967
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255967 557414 255978
rect 557470 255967 557538 256023
rect 557594 255967 557662 256023
rect 557718 255967 557786 256023
rect 557842 255978 597980 256023
rect 557842 255967 558474 255978
rect 528182 255922 558474 255967
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255899 597980 255922
rect -1916 255843 472732 255899
rect 472788 255843 472856 255899
rect 472912 255843 472980 255899
rect 473036 255843 473104 255899
rect 473160 255843 557414 255899
rect 557470 255843 557538 255899
rect 557594 255843 557662 255899
rect 557718 255843 557786 255899
rect 557842 255843 597980 255899
rect -1916 255826 597980 255843
rect 4156 248518 461204 248534
rect 4156 248462 4172 248518
rect 4228 248462 461132 248518
rect 461188 248462 461204 248518
rect 4156 248446 461204 248462
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 254994 244350
rect 255050 244294 255118 244350
rect 255174 244294 255242 244350
rect 255298 244294 255366 244350
rect 255422 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 361930 244350
rect 361986 244294 362054 244350
rect 362110 244294 362178 244350
rect 362234 244294 362302 244350
rect 362358 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 408594 244350
rect 408650 244294 408718 244350
rect 408774 244294 408842 244350
rect 408898 244294 408966 244350
rect 409022 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 446612 244350
rect 446668 244294 446736 244350
rect 446792 244294 446860 244350
rect 446916 244294 446984 244350
rect 447040 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 471932 244350
rect 471988 244294 472056 244350
rect 472112 244294 472180 244350
rect 472236 244294 472304 244350
rect 472360 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 556614 244350
rect 556670 244294 556738 244350
rect 556794 244294 556862 244350
rect 556918 244294 556986 244350
rect 557042 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 254994 244226
rect 255050 244170 255118 244226
rect 255174 244170 255242 244226
rect 255298 244170 255366 244226
rect 255422 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 361930 244226
rect 361986 244170 362054 244226
rect 362110 244170 362178 244226
rect 362234 244170 362302 244226
rect 362358 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 408594 244226
rect 408650 244170 408718 244226
rect 408774 244170 408842 244226
rect 408898 244170 408966 244226
rect 409022 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 446612 244226
rect 446668 244170 446736 244226
rect 446792 244170 446860 244226
rect 446916 244170 446984 244226
rect 447040 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 471932 244226
rect 471988 244170 472056 244226
rect 472112 244170 472180 244226
rect 472236 244170 472304 244226
rect 472360 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 556614 244226
rect 556670 244170 556738 244226
rect 556794 244170 556862 244226
rect 556918 244170 556986 244226
rect 557042 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 254994 244102
rect 255050 244046 255118 244102
rect 255174 244046 255242 244102
rect 255298 244046 255366 244102
rect 255422 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 361930 244102
rect 361986 244046 362054 244102
rect 362110 244046 362178 244102
rect 362234 244046 362302 244102
rect 362358 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 408594 244102
rect 408650 244046 408718 244102
rect 408774 244046 408842 244102
rect 408898 244046 408966 244102
rect 409022 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 446612 244102
rect 446668 244046 446736 244102
rect 446792 244046 446860 244102
rect 446916 244046 446984 244102
rect 447040 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 471932 244102
rect 471988 244046 472056 244102
rect 472112 244046 472180 244102
rect 472236 244046 472304 244102
rect 472360 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 556614 244102
rect 556670 244046 556738 244102
rect 556794 244046 556862 244102
rect 556918 244046 556986 244102
rect 557042 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 254994 243978
rect 255050 243922 255118 243978
rect 255174 243922 255242 243978
rect 255298 243922 255366 243978
rect 255422 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 361930 243978
rect 361986 243922 362054 243978
rect 362110 243922 362178 243978
rect 362234 243922 362302 243978
rect 362358 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 408594 243978
rect 408650 243922 408718 243978
rect 408774 243922 408842 243978
rect 408898 243922 408966 243978
rect 409022 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 446612 243978
rect 446668 243922 446736 243978
rect 446792 243922 446860 243978
rect 446916 243922 446984 243978
rect 447040 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 471932 243978
rect 471988 243922 472056 243978
rect 472112 243922 472180 243978
rect 472236 243922 472304 243978
rect 472360 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 556614 243978
rect 556670 243922 556738 243978
rect 556794 243922 556862 243978
rect 556918 243922 556986 243978
rect 557042 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 361130 238350
rect 361186 238294 361254 238350
rect 361310 238294 361378 238350
rect 361434 238294 361502 238350
rect 361558 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 404874 238350
rect 404930 238294 404998 238350
rect 405054 238294 405122 238350
rect 405178 238294 405246 238350
rect 405302 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 445812 238350
rect 445868 238294 445936 238350
rect 445992 238294 446060 238350
rect 446116 238294 446184 238350
rect 446240 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 472732 238350
rect 472788 238294 472856 238350
rect 472912 238294 472980 238350
rect 473036 238294 473104 238350
rect 473160 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 557414 238350
rect 557470 238294 557538 238350
rect 557594 238294 557662 238350
rect 557718 238294 557786 238350
rect 557842 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 361130 238226
rect 361186 238170 361254 238226
rect 361310 238170 361378 238226
rect 361434 238170 361502 238226
rect 361558 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 404874 238226
rect 404930 238170 404998 238226
rect 405054 238170 405122 238226
rect 405178 238170 405246 238226
rect 405302 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 445812 238226
rect 445868 238170 445936 238226
rect 445992 238170 446060 238226
rect 446116 238170 446184 238226
rect 446240 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 472732 238226
rect 472788 238170 472856 238226
rect 472912 238170 472980 238226
rect 473036 238170 473104 238226
rect 473160 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 557414 238226
rect 557470 238170 557538 238226
rect 557594 238170 557662 238226
rect 557718 238170 557786 238226
rect 557842 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 361130 238102
rect 361186 238046 361254 238102
rect 361310 238046 361378 238102
rect 361434 238046 361502 238102
rect 361558 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 404874 238102
rect 404930 238046 404998 238102
rect 405054 238046 405122 238102
rect 405178 238046 405246 238102
rect 405302 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 445812 238102
rect 445868 238046 445936 238102
rect 445992 238046 446060 238102
rect 446116 238046 446184 238102
rect 446240 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 472732 238102
rect 472788 238046 472856 238102
rect 472912 238046 472980 238102
rect 473036 238046 473104 238102
rect 473160 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 557414 238102
rect 557470 238046 557538 238102
rect 557594 238046 557662 238102
rect 557718 238046 557786 238102
rect 557842 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 361130 237978
rect 361186 237922 361254 237978
rect 361310 237922 361378 237978
rect 361434 237922 361502 237978
rect 361558 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 404874 237978
rect 404930 237922 404998 237978
rect 405054 237922 405122 237978
rect 405178 237922 405246 237978
rect 405302 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 445812 237978
rect 445868 237922 445936 237978
rect 445992 237922 446060 237978
rect 446116 237922 446184 237978
rect 446240 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 472732 237978
rect 472788 237922 472856 237978
rect 472912 237922 472980 237978
rect 473036 237922 473104 237978
rect 473160 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 557414 237978
rect 557470 237922 557538 237978
rect 557594 237922 557662 237978
rect 557718 237922 557786 237978
rect 557842 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect 4156 235198 464676 235214
rect 4156 235142 4172 235198
rect 4228 235142 464604 235198
rect 464660 235142 464676 235198
rect 4156 235126 464676 235142
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 361930 226350
rect 361986 226294 362054 226350
rect 362110 226294 362178 226350
rect 362234 226294 362302 226350
rect 362358 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 408594 226350
rect 408650 226294 408718 226350
rect 408774 226294 408842 226350
rect 408898 226294 408966 226350
rect 409022 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 446612 226350
rect 446668 226294 446736 226350
rect 446792 226294 446860 226350
rect 446916 226294 446984 226350
rect 447040 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 471932 226350
rect 471988 226294 472056 226350
rect 472112 226294 472180 226350
rect 472236 226294 472304 226350
rect 472360 226294 500754 226350
rect 500810 226294 500878 226350
rect 500934 226294 501002 226350
rect 501058 226294 501126 226350
rect 501182 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 556614 226350
rect 556670 226294 556738 226350
rect 556794 226294 556862 226350
rect 556918 226294 556986 226350
rect 557042 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 361930 226226
rect 361986 226170 362054 226226
rect 362110 226170 362178 226226
rect 362234 226170 362302 226226
rect 362358 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 408594 226226
rect 408650 226170 408718 226226
rect 408774 226170 408842 226226
rect 408898 226170 408966 226226
rect 409022 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 446612 226226
rect 446668 226170 446736 226226
rect 446792 226170 446860 226226
rect 446916 226170 446984 226226
rect 447040 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 471932 226226
rect 471988 226170 472056 226226
rect 472112 226170 472180 226226
rect 472236 226170 472304 226226
rect 472360 226170 500754 226226
rect 500810 226170 500878 226226
rect 500934 226170 501002 226226
rect 501058 226170 501126 226226
rect 501182 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 556614 226226
rect 556670 226170 556738 226226
rect 556794 226170 556862 226226
rect 556918 226170 556986 226226
rect 557042 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 361930 226102
rect 361986 226046 362054 226102
rect 362110 226046 362178 226102
rect 362234 226046 362302 226102
rect 362358 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 408594 226102
rect 408650 226046 408718 226102
rect 408774 226046 408842 226102
rect 408898 226046 408966 226102
rect 409022 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 446612 226102
rect 446668 226046 446736 226102
rect 446792 226046 446860 226102
rect 446916 226046 446984 226102
rect 447040 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 471932 226102
rect 471988 226046 472056 226102
rect 472112 226046 472180 226102
rect 472236 226046 472304 226102
rect 472360 226046 500754 226102
rect 500810 226046 500878 226102
rect 500934 226046 501002 226102
rect 501058 226046 501126 226102
rect 501182 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 556614 226102
rect 556670 226046 556738 226102
rect 556794 226046 556862 226102
rect 556918 226046 556986 226102
rect 557042 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 361930 225978
rect 361986 225922 362054 225978
rect 362110 225922 362178 225978
rect 362234 225922 362302 225978
rect 362358 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 408594 225978
rect 408650 225922 408718 225978
rect 408774 225922 408842 225978
rect 408898 225922 408966 225978
rect 409022 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 446612 225978
rect 446668 225922 446736 225978
rect 446792 225922 446860 225978
rect 446916 225922 446984 225978
rect 447040 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 471932 225978
rect 471988 225922 472056 225978
rect 472112 225922 472180 225978
rect 472236 225922 472304 225978
rect 472360 225922 500754 225978
rect 500810 225922 500878 225978
rect 500934 225922 501002 225978
rect 501058 225922 501126 225978
rect 501182 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 556614 225978
rect 556670 225922 556738 225978
rect 556794 225922 556862 225978
rect 556918 225922 556986 225978
rect 557042 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 361130 220350
rect 361186 220294 361254 220350
rect 361310 220294 361378 220350
rect 361434 220294 361502 220350
rect 361558 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 404874 220350
rect 404930 220294 404998 220350
rect 405054 220294 405122 220350
rect 405178 220294 405246 220350
rect 405302 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 445812 220350
rect 445868 220294 445936 220350
rect 445992 220294 446060 220350
rect 446116 220294 446184 220350
rect 446240 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 472732 220350
rect 472788 220294 472856 220350
rect 472912 220294 472980 220350
rect 473036 220294 473104 220350
rect 473160 220294 497034 220350
rect 497090 220294 497158 220350
rect 497214 220294 497282 220350
rect 497338 220294 497406 220350
rect 497462 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 557414 220350
rect 557470 220294 557538 220350
rect 557594 220294 557662 220350
rect 557718 220294 557786 220350
rect 557842 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 361130 220226
rect 361186 220170 361254 220226
rect 361310 220170 361378 220226
rect 361434 220170 361502 220226
rect 361558 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 404874 220226
rect 404930 220170 404998 220226
rect 405054 220170 405122 220226
rect 405178 220170 405246 220226
rect 405302 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 445812 220226
rect 445868 220170 445936 220226
rect 445992 220170 446060 220226
rect 446116 220170 446184 220226
rect 446240 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 472732 220226
rect 472788 220170 472856 220226
rect 472912 220170 472980 220226
rect 473036 220170 473104 220226
rect 473160 220170 497034 220226
rect 497090 220170 497158 220226
rect 497214 220170 497282 220226
rect 497338 220170 497406 220226
rect 497462 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 557414 220226
rect 557470 220170 557538 220226
rect 557594 220170 557662 220226
rect 557718 220170 557786 220226
rect 557842 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 361130 220102
rect 361186 220046 361254 220102
rect 361310 220046 361378 220102
rect 361434 220046 361502 220102
rect 361558 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 404874 220102
rect 404930 220046 404998 220102
rect 405054 220046 405122 220102
rect 405178 220046 405246 220102
rect 405302 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 445812 220102
rect 445868 220046 445936 220102
rect 445992 220046 446060 220102
rect 446116 220046 446184 220102
rect 446240 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 472732 220102
rect 472788 220046 472856 220102
rect 472912 220046 472980 220102
rect 473036 220046 473104 220102
rect 473160 220046 497034 220102
rect 497090 220046 497158 220102
rect 497214 220046 497282 220102
rect 497338 220046 497406 220102
rect 497462 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 557414 220102
rect 557470 220046 557538 220102
rect 557594 220046 557662 220102
rect 557718 220046 557786 220102
rect 557842 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 361130 219978
rect 361186 219922 361254 219978
rect 361310 219922 361378 219978
rect 361434 219922 361502 219978
rect 361558 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 404874 219978
rect 404930 219922 404998 219978
rect 405054 219922 405122 219978
rect 405178 219922 405246 219978
rect 405302 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 445812 219978
rect 445868 219922 445936 219978
rect 445992 219922 446060 219978
rect 446116 219922 446184 219978
rect 446240 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 472732 219978
rect 472788 219922 472856 219978
rect 472912 219922 472980 219978
rect 473036 219922 473104 219978
rect 473160 219922 497034 219978
rect 497090 219922 497158 219978
rect 497214 219922 497282 219978
rect 497338 219922 497406 219978
rect 497462 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 557414 219978
rect 557470 219922 557538 219978
rect 557594 219922 557662 219978
rect 557718 219922 557786 219978
rect 557842 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 101394 208350
rect 101450 208294 101518 208350
rect 101574 208294 101642 208350
rect 101698 208294 101766 208350
rect 101822 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 224274 208350
rect 224330 208294 224398 208350
rect 224454 208294 224522 208350
rect 224578 208294 224646 208350
rect 224702 208294 254994 208350
rect 255050 208294 255118 208350
rect 255174 208294 255242 208350
rect 255298 208294 255366 208350
rect 255422 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 361930 208350
rect 361986 208294 362054 208350
rect 362110 208294 362178 208350
rect 362234 208294 362302 208350
rect 362358 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208294 408594 208350
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 446612 208350
rect 446668 208294 446736 208350
rect 446792 208294 446860 208350
rect 446916 208294 446984 208350
rect 447040 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 471932 208350
rect 471988 208294 472056 208350
rect 472112 208294 472180 208350
rect 472236 208294 472304 208350
rect 472360 208294 500754 208350
rect 500810 208294 500878 208350
rect 500934 208294 501002 208350
rect 501058 208294 501126 208350
rect 501182 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 556614 208350
rect 556670 208294 556738 208350
rect 556794 208294 556862 208350
rect 556918 208294 556986 208350
rect 557042 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 101394 208226
rect 101450 208170 101518 208226
rect 101574 208170 101642 208226
rect 101698 208170 101766 208226
rect 101822 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 224274 208226
rect 224330 208170 224398 208226
rect 224454 208170 224522 208226
rect 224578 208170 224646 208226
rect 224702 208170 254994 208226
rect 255050 208170 255118 208226
rect 255174 208170 255242 208226
rect 255298 208170 255366 208226
rect 255422 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 361930 208226
rect 361986 208170 362054 208226
rect 362110 208170 362178 208226
rect 362234 208170 362302 208226
rect 362358 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208170 408594 208226
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 446612 208226
rect 446668 208170 446736 208226
rect 446792 208170 446860 208226
rect 446916 208170 446984 208226
rect 447040 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 471932 208226
rect 471988 208170 472056 208226
rect 472112 208170 472180 208226
rect 472236 208170 472304 208226
rect 472360 208170 500754 208226
rect 500810 208170 500878 208226
rect 500934 208170 501002 208226
rect 501058 208170 501126 208226
rect 501182 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 556614 208226
rect 556670 208170 556738 208226
rect 556794 208170 556862 208226
rect 556918 208170 556986 208226
rect 557042 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 101394 208102
rect 101450 208046 101518 208102
rect 101574 208046 101642 208102
rect 101698 208046 101766 208102
rect 101822 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 224274 208102
rect 224330 208046 224398 208102
rect 224454 208046 224522 208102
rect 224578 208046 224646 208102
rect 224702 208046 254994 208102
rect 255050 208046 255118 208102
rect 255174 208046 255242 208102
rect 255298 208046 255366 208102
rect 255422 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 361930 208102
rect 361986 208046 362054 208102
rect 362110 208046 362178 208102
rect 362234 208046 362302 208102
rect 362358 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 446612 208102
rect 446668 208046 446736 208102
rect 446792 208046 446860 208102
rect 446916 208046 446984 208102
rect 447040 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 471932 208102
rect 471988 208046 472056 208102
rect 472112 208046 472180 208102
rect 472236 208046 472304 208102
rect 472360 208046 500754 208102
rect 500810 208046 500878 208102
rect 500934 208046 501002 208102
rect 501058 208046 501126 208102
rect 501182 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 556614 208102
rect 556670 208046 556738 208102
rect 556794 208046 556862 208102
rect 556918 208046 556986 208102
rect 557042 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 101394 207978
rect 101450 207922 101518 207978
rect 101574 207922 101642 207978
rect 101698 207922 101766 207978
rect 101822 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 224274 207978
rect 224330 207922 224398 207978
rect 224454 207922 224522 207978
rect 224578 207922 224646 207978
rect 224702 207922 254994 207978
rect 255050 207922 255118 207978
rect 255174 207922 255242 207978
rect 255298 207922 255366 207978
rect 255422 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 361930 207978
rect 361986 207922 362054 207978
rect 362110 207922 362178 207978
rect 362234 207922 362302 207978
rect 362358 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 446612 207978
rect 446668 207922 446736 207978
rect 446792 207922 446860 207978
rect 446916 207922 446984 207978
rect 447040 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 471932 207978
rect 471988 207922 472056 207978
rect 472112 207922 472180 207978
rect 472236 207922 472304 207978
rect 472360 207922 500754 207978
rect 500810 207922 500878 207978
rect 500934 207922 501002 207978
rect 501058 207922 501126 207978
rect 501182 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 556614 207978
rect 556670 207922 556738 207978
rect 556794 207922 556862 207978
rect 556918 207922 556986 207978
rect 557042 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect 4156 206578 464564 206594
rect 4156 206522 4172 206578
rect 4228 206522 464492 206578
rect 464548 206522 464564 206578
rect 4156 206506 464564 206522
rect 284828 206398 590228 206414
rect 284828 206342 284844 206398
rect 284900 206342 590156 206398
rect 590212 206342 590228 206398
rect 284828 206326 590228 206342
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 64518 202350
rect 64574 202294 64642 202350
rect 64698 202294 66954 202350
rect 67010 202294 67078 202350
rect 67134 202294 67202 202350
rect 67258 202294 67326 202350
rect 67382 202294 95238 202350
rect 95294 202294 95362 202350
rect 95418 202294 97674 202350
rect 97730 202294 97798 202350
rect 97854 202294 97922 202350
rect 97978 202294 98046 202350
rect 98102 202294 125958 202350
rect 126014 202294 126082 202350
rect 126138 202294 128394 202350
rect 128450 202294 128518 202350
rect 128574 202294 128642 202350
rect 128698 202294 128766 202350
rect 128822 202294 156678 202350
rect 156734 202294 156802 202350
rect 156858 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 187398 202350
rect 187454 202294 187522 202350
rect 187578 202294 189834 202350
rect 189890 202294 189958 202350
rect 190014 202294 190082 202350
rect 190138 202294 190206 202350
rect 190262 202294 218118 202350
rect 218174 202294 218242 202350
rect 218298 202294 220554 202350
rect 220610 202294 220678 202350
rect 220734 202294 220802 202350
rect 220858 202294 220926 202350
rect 220982 202294 248838 202350
rect 248894 202294 248962 202350
rect 249018 202294 251274 202350
rect 251330 202294 251398 202350
rect 251454 202294 251522 202350
rect 251578 202294 251646 202350
rect 251702 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 361130 202350
rect 361186 202294 361254 202350
rect 361310 202294 361378 202350
rect 361434 202294 361502 202350
rect 361558 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 445812 202350
rect 445868 202294 445936 202350
rect 445992 202294 446060 202350
rect 446116 202294 446184 202350
rect 446240 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 472732 202350
rect 472788 202294 472856 202350
rect 472912 202294 472980 202350
rect 473036 202294 473104 202350
rect 473160 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 557414 202350
rect 557470 202294 557538 202350
rect 557594 202294 557662 202350
rect 557718 202294 557786 202350
rect 557842 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 64518 202226
rect 64574 202170 64642 202226
rect 64698 202170 66954 202226
rect 67010 202170 67078 202226
rect 67134 202170 67202 202226
rect 67258 202170 67326 202226
rect 67382 202170 95238 202226
rect 95294 202170 95362 202226
rect 95418 202170 97674 202226
rect 97730 202170 97798 202226
rect 97854 202170 97922 202226
rect 97978 202170 98046 202226
rect 98102 202170 125958 202226
rect 126014 202170 126082 202226
rect 126138 202170 128394 202226
rect 128450 202170 128518 202226
rect 128574 202170 128642 202226
rect 128698 202170 128766 202226
rect 128822 202170 156678 202226
rect 156734 202170 156802 202226
rect 156858 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 187398 202226
rect 187454 202170 187522 202226
rect 187578 202170 189834 202226
rect 189890 202170 189958 202226
rect 190014 202170 190082 202226
rect 190138 202170 190206 202226
rect 190262 202170 218118 202226
rect 218174 202170 218242 202226
rect 218298 202170 220554 202226
rect 220610 202170 220678 202226
rect 220734 202170 220802 202226
rect 220858 202170 220926 202226
rect 220982 202170 248838 202226
rect 248894 202170 248962 202226
rect 249018 202170 251274 202226
rect 251330 202170 251398 202226
rect 251454 202170 251522 202226
rect 251578 202170 251646 202226
rect 251702 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 361130 202226
rect 361186 202170 361254 202226
rect 361310 202170 361378 202226
rect 361434 202170 361502 202226
rect 361558 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 445812 202226
rect 445868 202170 445936 202226
rect 445992 202170 446060 202226
rect 446116 202170 446184 202226
rect 446240 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 472732 202226
rect 472788 202170 472856 202226
rect 472912 202170 472980 202226
rect 473036 202170 473104 202226
rect 473160 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 557414 202226
rect 557470 202170 557538 202226
rect 557594 202170 557662 202226
rect 557718 202170 557786 202226
rect 557842 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 64518 202102
rect 64574 202046 64642 202102
rect 64698 202046 66954 202102
rect 67010 202046 67078 202102
rect 67134 202046 67202 202102
rect 67258 202046 67326 202102
rect 67382 202046 95238 202102
rect 95294 202046 95362 202102
rect 95418 202046 97674 202102
rect 97730 202046 97798 202102
rect 97854 202046 97922 202102
rect 97978 202046 98046 202102
rect 98102 202046 125958 202102
rect 126014 202046 126082 202102
rect 126138 202046 128394 202102
rect 128450 202046 128518 202102
rect 128574 202046 128642 202102
rect 128698 202046 128766 202102
rect 128822 202046 156678 202102
rect 156734 202046 156802 202102
rect 156858 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 187398 202102
rect 187454 202046 187522 202102
rect 187578 202046 189834 202102
rect 189890 202046 189958 202102
rect 190014 202046 190082 202102
rect 190138 202046 190206 202102
rect 190262 202046 218118 202102
rect 218174 202046 218242 202102
rect 218298 202046 220554 202102
rect 220610 202046 220678 202102
rect 220734 202046 220802 202102
rect 220858 202046 220926 202102
rect 220982 202046 248838 202102
rect 248894 202046 248962 202102
rect 249018 202046 251274 202102
rect 251330 202046 251398 202102
rect 251454 202046 251522 202102
rect 251578 202046 251646 202102
rect 251702 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 361130 202102
rect 361186 202046 361254 202102
rect 361310 202046 361378 202102
rect 361434 202046 361502 202102
rect 361558 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 445812 202102
rect 445868 202046 445936 202102
rect 445992 202046 446060 202102
rect 446116 202046 446184 202102
rect 446240 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 472732 202102
rect 472788 202046 472856 202102
rect 472912 202046 472980 202102
rect 473036 202046 473104 202102
rect 473160 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 557414 202102
rect 557470 202046 557538 202102
rect 557594 202046 557662 202102
rect 557718 202046 557786 202102
rect 557842 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 64518 201978
rect 64574 201922 64642 201978
rect 64698 201922 66954 201978
rect 67010 201922 67078 201978
rect 67134 201922 67202 201978
rect 67258 201922 67326 201978
rect 67382 201922 95238 201978
rect 95294 201922 95362 201978
rect 95418 201922 97674 201978
rect 97730 201922 97798 201978
rect 97854 201922 97922 201978
rect 97978 201922 98046 201978
rect 98102 201922 125958 201978
rect 126014 201922 126082 201978
rect 126138 201922 128394 201978
rect 128450 201922 128518 201978
rect 128574 201922 128642 201978
rect 128698 201922 128766 201978
rect 128822 201922 156678 201978
rect 156734 201922 156802 201978
rect 156858 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 187398 201978
rect 187454 201922 187522 201978
rect 187578 201922 189834 201978
rect 189890 201922 189958 201978
rect 190014 201922 190082 201978
rect 190138 201922 190206 201978
rect 190262 201922 218118 201978
rect 218174 201922 218242 201978
rect 218298 201922 220554 201978
rect 220610 201922 220678 201978
rect 220734 201922 220802 201978
rect 220858 201922 220926 201978
rect 220982 201922 248838 201978
rect 248894 201922 248962 201978
rect 249018 201922 251274 201978
rect 251330 201922 251398 201978
rect 251454 201922 251522 201978
rect 251578 201922 251646 201978
rect 251702 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 361130 201978
rect 361186 201922 361254 201978
rect 361310 201922 361378 201978
rect 361434 201922 361502 201978
rect 361558 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 445812 201978
rect 445868 201922 445936 201978
rect 445992 201922 446060 201978
rect 446116 201922 446184 201978
rect 446240 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 472732 201978
rect 472788 201922 472856 201978
rect 472912 201922 472980 201978
rect 473036 201922 473104 201978
rect 473160 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 557414 201978
rect 557470 201922 557538 201978
rect 557594 201922 557662 201978
rect 557718 201922 557786 201978
rect 557842 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 70674 190350
rect 70730 190294 70798 190350
rect 70854 190294 70922 190350
rect 70978 190294 71046 190350
rect 71102 190294 79878 190350
rect 79934 190294 80002 190350
rect 80058 190294 101394 190350
rect 101450 190294 101518 190350
rect 101574 190294 101642 190350
rect 101698 190294 101766 190350
rect 101822 190294 110598 190350
rect 110654 190294 110722 190350
rect 110778 190294 132114 190350
rect 132170 190294 132238 190350
rect 132294 190294 132362 190350
rect 132418 190294 132486 190350
rect 132542 190294 141318 190350
rect 141374 190294 141442 190350
rect 141498 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 172038 190350
rect 172094 190294 172162 190350
rect 172218 190294 193554 190350
rect 193610 190294 193678 190350
rect 193734 190294 193802 190350
rect 193858 190294 193926 190350
rect 193982 190294 202758 190350
rect 202814 190294 202882 190350
rect 202938 190294 224274 190350
rect 224330 190294 224398 190350
rect 224454 190294 224522 190350
rect 224578 190294 224646 190350
rect 224702 190294 233478 190350
rect 233534 190294 233602 190350
rect 233658 190294 254994 190350
rect 255050 190294 255118 190350
rect 255174 190294 255242 190350
rect 255298 190294 255366 190350
rect 255422 190294 264198 190350
rect 264254 190294 264322 190350
rect 264378 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 361930 190350
rect 361986 190294 362054 190350
rect 362110 190294 362178 190350
rect 362234 190294 362302 190350
rect 362358 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 446612 190350
rect 446668 190294 446736 190350
rect 446792 190294 446860 190350
rect 446916 190294 446984 190350
rect 447040 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 471932 190350
rect 471988 190294 472056 190350
rect 472112 190294 472180 190350
rect 472236 190294 472304 190350
rect 472360 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 556614 190350
rect 556670 190294 556738 190350
rect 556794 190294 556862 190350
rect 556918 190294 556986 190350
rect 557042 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 70674 190226
rect 70730 190170 70798 190226
rect 70854 190170 70922 190226
rect 70978 190170 71046 190226
rect 71102 190170 79878 190226
rect 79934 190170 80002 190226
rect 80058 190170 101394 190226
rect 101450 190170 101518 190226
rect 101574 190170 101642 190226
rect 101698 190170 101766 190226
rect 101822 190170 110598 190226
rect 110654 190170 110722 190226
rect 110778 190170 132114 190226
rect 132170 190170 132238 190226
rect 132294 190170 132362 190226
rect 132418 190170 132486 190226
rect 132542 190170 141318 190226
rect 141374 190170 141442 190226
rect 141498 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 172038 190226
rect 172094 190170 172162 190226
rect 172218 190170 193554 190226
rect 193610 190170 193678 190226
rect 193734 190170 193802 190226
rect 193858 190170 193926 190226
rect 193982 190170 202758 190226
rect 202814 190170 202882 190226
rect 202938 190170 224274 190226
rect 224330 190170 224398 190226
rect 224454 190170 224522 190226
rect 224578 190170 224646 190226
rect 224702 190170 233478 190226
rect 233534 190170 233602 190226
rect 233658 190170 254994 190226
rect 255050 190170 255118 190226
rect 255174 190170 255242 190226
rect 255298 190170 255366 190226
rect 255422 190170 264198 190226
rect 264254 190170 264322 190226
rect 264378 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 361930 190226
rect 361986 190170 362054 190226
rect 362110 190170 362178 190226
rect 362234 190170 362302 190226
rect 362358 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 446612 190226
rect 446668 190170 446736 190226
rect 446792 190170 446860 190226
rect 446916 190170 446984 190226
rect 447040 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 471932 190226
rect 471988 190170 472056 190226
rect 472112 190170 472180 190226
rect 472236 190170 472304 190226
rect 472360 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 556614 190226
rect 556670 190170 556738 190226
rect 556794 190170 556862 190226
rect 556918 190170 556986 190226
rect 557042 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 70674 190102
rect 70730 190046 70798 190102
rect 70854 190046 70922 190102
rect 70978 190046 71046 190102
rect 71102 190046 79878 190102
rect 79934 190046 80002 190102
rect 80058 190046 101394 190102
rect 101450 190046 101518 190102
rect 101574 190046 101642 190102
rect 101698 190046 101766 190102
rect 101822 190046 110598 190102
rect 110654 190046 110722 190102
rect 110778 190046 132114 190102
rect 132170 190046 132238 190102
rect 132294 190046 132362 190102
rect 132418 190046 132486 190102
rect 132542 190046 141318 190102
rect 141374 190046 141442 190102
rect 141498 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 172038 190102
rect 172094 190046 172162 190102
rect 172218 190046 193554 190102
rect 193610 190046 193678 190102
rect 193734 190046 193802 190102
rect 193858 190046 193926 190102
rect 193982 190046 202758 190102
rect 202814 190046 202882 190102
rect 202938 190046 224274 190102
rect 224330 190046 224398 190102
rect 224454 190046 224522 190102
rect 224578 190046 224646 190102
rect 224702 190046 233478 190102
rect 233534 190046 233602 190102
rect 233658 190046 254994 190102
rect 255050 190046 255118 190102
rect 255174 190046 255242 190102
rect 255298 190046 255366 190102
rect 255422 190046 264198 190102
rect 264254 190046 264322 190102
rect 264378 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 361930 190102
rect 361986 190046 362054 190102
rect 362110 190046 362178 190102
rect 362234 190046 362302 190102
rect 362358 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 446612 190102
rect 446668 190046 446736 190102
rect 446792 190046 446860 190102
rect 446916 190046 446984 190102
rect 447040 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 471932 190102
rect 471988 190046 472056 190102
rect 472112 190046 472180 190102
rect 472236 190046 472304 190102
rect 472360 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 556614 190102
rect 556670 190046 556738 190102
rect 556794 190046 556862 190102
rect 556918 190046 556986 190102
rect 557042 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 70674 189978
rect 70730 189922 70798 189978
rect 70854 189922 70922 189978
rect 70978 189922 71046 189978
rect 71102 189922 79878 189978
rect 79934 189922 80002 189978
rect 80058 189922 101394 189978
rect 101450 189922 101518 189978
rect 101574 189922 101642 189978
rect 101698 189922 101766 189978
rect 101822 189922 110598 189978
rect 110654 189922 110722 189978
rect 110778 189922 132114 189978
rect 132170 189922 132238 189978
rect 132294 189922 132362 189978
rect 132418 189922 132486 189978
rect 132542 189922 141318 189978
rect 141374 189922 141442 189978
rect 141498 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 172038 189978
rect 172094 189922 172162 189978
rect 172218 189922 193554 189978
rect 193610 189922 193678 189978
rect 193734 189922 193802 189978
rect 193858 189922 193926 189978
rect 193982 189922 202758 189978
rect 202814 189922 202882 189978
rect 202938 189922 224274 189978
rect 224330 189922 224398 189978
rect 224454 189922 224522 189978
rect 224578 189922 224646 189978
rect 224702 189922 233478 189978
rect 233534 189922 233602 189978
rect 233658 189922 254994 189978
rect 255050 189922 255118 189978
rect 255174 189922 255242 189978
rect 255298 189922 255366 189978
rect 255422 189922 264198 189978
rect 264254 189922 264322 189978
rect 264378 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 361930 189978
rect 361986 189922 362054 189978
rect 362110 189922 362178 189978
rect 362234 189922 362302 189978
rect 362358 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 446612 189978
rect 446668 189922 446736 189978
rect 446792 189922 446860 189978
rect 446916 189922 446984 189978
rect 447040 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 471932 189978
rect 471988 189922 472056 189978
rect 472112 189922 472180 189978
rect 472236 189922 472304 189978
rect 472360 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 556614 189978
rect 556670 189922 556738 189978
rect 556794 189922 556862 189978
rect 556918 189922 556986 189978
rect 557042 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 64518 184350
rect 64574 184294 64642 184350
rect 64698 184294 66954 184350
rect 67010 184294 67078 184350
rect 67134 184294 67202 184350
rect 67258 184294 67326 184350
rect 67382 184294 95238 184350
rect 95294 184294 95362 184350
rect 95418 184294 97674 184350
rect 97730 184294 97798 184350
rect 97854 184294 97922 184350
rect 97978 184294 98046 184350
rect 98102 184294 125958 184350
rect 126014 184294 126082 184350
rect 126138 184294 128394 184350
rect 128450 184294 128518 184350
rect 128574 184294 128642 184350
rect 128698 184294 128766 184350
rect 128822 184294 156678 184350
rect 156734 184294 156802 184350
rect 156858 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 187398 184350
rect 187454 184294 187522 184350
rect 187578 184294 189834 184350
rect 189890 184294 189958 184350
rect 190014 184294 190082 184350
rect 190138 184294 190206 184350
rect 190262 184294 218118 184350
rect 218174 184294 218242 184350
rect 218298 184294 220554 184350
rect 220610 184294 220678 184350
rect 220734 184294 220802 184350
rect 220858 184294 220926 184350
rect 220982 184294 248838 184350
rect 248894 184294 248962 184350
rect 249018 184294 251274 184350
rect 251330 184294 251398 184350
rect 251454 184294 251522 184350
rect 251578 184294 251646 184350
rect 251702 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 361130 184350
rect 361186 184294 361254 184350
rect 361310 184294 361378 184350
rect 361434 184294 361502 184350
rect 361558 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 404874 184350
rect 404930 184294 404998 184350
rect 405054 184294 405122 184350
rect 405178 184294 405246 184350
rect 405302 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 445812 184350
rect 445868 184294 445936 184350
rect 445992 184294 446060 184350
rect 446116 184294 446184 184350
rect 446240 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 472732 184350
rect 472788 184294 472856 184350
rect 472912 184294 472980 184350
rect 473036 184294 473104 184350
rect 473160 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 557414 184350
rect 557470 184294 557538 184350
rect 557594 184294 557662 184350
rect 557718 184294 557786 184350
rect 557842 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 64518 184226
rect 64574 184170 64642 184226
rect 64698 184170 66954 184226
rect 67010 184170 67078 184226
rect 67134 184170 67202 184226
rect 67258 184170 67326 184226
rect 67382 184170 95238 184226
rect 95294 184170 95362 184226
rect 95418 184170 97674 184226
rect 97730 184170 97798 184226
rect 97854 184170 97922 184226
rect 97978 184170 98046 184226
rect 98102 184170 125958 184226
rect 126014 184170 126082 184226
rect 126138 184170 128394 184226
rect 128450 184170 128518 184226
rect 128574 184170 128642 184226
rect 128698 184170 128766 184226
rect 128822 184170 156678 184226
rect 156734 184170 156802 184226
rect 156858 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 187398 184226
rect 187454 184170 187522 184226
rect 187578 184170 189834 184226
rect 189890 184170 189958 184226
rect 190014 184170 190082 184226
rect 190138 184170 190206 184226
rect 190262 184170 218118 184226
rect 218174 184170 218242 184226
rect 218298 184170 220554 184226
rect 220610 184170 220678 184226
rect 220734 184170 220802 184226
rect 220858 184170 220926 184226
rect 220982 184170 248838 184226
rect 248894 184170 248962 184226
rect 249018 184170 251274 184226
rect 251330 184170 251398 184226
rect 251454 184170 251522 184226
rect 251578 184170 251646 184226
rect 251702 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 361130 184226
rect 361186 184170 361254 184226
rect 361310 184170 361378 184226
rect 361434 184170 361502 184226
rect 361558 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 404874 184226
rect 404930 184170 404998 184226
rect 405054 184170 405122 184226
rect 405178 184170 405246 184226
rect 405302 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 445812 184226
rect 445868 184170 445936 184226
rect 445992 184170 446060 184226
rect 446116 184170 446184 184226
rect 446240 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 472732 184226
rect 472788 184170 472856 184226
rect 472912 184170 472980 184226
rect 473036 184170 473104 184226
rect 473160 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 557414 184226
rect 557470 184170 557538 184226
rect 557594 184170 557662 184226
rect 557718 184170 557786 184226
rect 557842 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 64518 184102
rect 64574 184046 64642 184102
rect 64698 184046 66954 184102
rect 67010 184046 67078 184102
rect 67134 184046 67202 184102
rect 67258 184046 67326 184102
rect 67382 184046 95238 184102
rect 95294 184046 95362 184102
rect 95418 184046 97674 184102
rect 97730 184046 97798 184102
rect 97854 184046 97922 184102
rect 97978 184046 98046 184102
rect 98102 184046 125958 184102
rect 126014 184046 126082 184102
rect 126138 184046 128394 184102
rect 128450 184046 128518 184102
rect 128574 184046 128642 184102
rect 128698 184046 128766 184102
rect 128822 184046 156678 184102
rect 156734 184046 156802 184102
rect 156858 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 187398 184102
rect 187454 184046 187522 184102
rect 187578 184046 189834 184102
rect 189890 184046 189958 184102
rect 190014 184046 190082 184102
rect 190138 184046 190206 184102
rect 190262 184046 218118 184102
rect 218174 184046 218242 184102
rect 218298 184046 220554 184102
rect 220610 184046 220678 184102
rect 220734 184046 220802 184102
rect 220858 184046 220926 184102
rect 220982 184046 248838 184102
rect 248894 184046 248962 184102
rect 249018 184046 251274 184102
rect 251330 184046 251398 184102
rect 251454 184046 251522 184102
rect 251578 184046 251646 184102
rect 251702 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 361130 184102
rect 361186 184046 361254 184102
rect 361310 184046 361378 184102
rect 361434 184046 361502 184102
rect 361558 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 404874 184102
rect 404930 184046 404998 184102
rect 405054 184046 405122 184102
rect 405178 184046 405246 184102
rect 405302 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 445812 184102
rect 445868 184046 445936 184102
rect 445992 184046 446060 184102
rect 446116 184046 446184 184102
rect 446240 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 472732 184102
rect 472788 184046 472856 184102
rect 472912 184046 472980 184102
rect 473036 184046 473104 184102
rect 473160 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 557414 184102
rect 557470 184046 557538 184102
rect 557594 184046 557662 184102
rect 557718 184046 557786 184102
rect 557842 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 64518 183978
rect 64574 183922 64642 183978
rect 64698 183922 66954 183978
rect 67010 183922 67078 183978
rect 67134 183922 67202 183978
rect 67258 183922 67326 183978
rect 67382 183922 95238 183978
rect 95294 183922 95362 183978
rect 95418 183922 97674 183978
rect 97730 183922 97798 183978
rect 97854 183922 97922 183978
rect 97978 183922 98046 183978
rect 98102 183922 125958 183978
rect 126014 183922 126082 183978
rect 126138 183922 128394 183978
rect 128450 183922 128518 183978
rect 128574 183922 128642 183978
rect 128698 183922 128766 183978
rect 128822 183922 156678 183978
rect 156734 183922 156802 183978
rect 156858 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 187398 183978
rect 187454 183922 187522 183978
rect 187578 183922 189834 183978
rect 189890 183922 189958 183978
rect 190014 183922 190082 183978
rect 190138 183922 190206 183978
rect 190262 183922 218118 183978
rect 218174 183922 218242 183978
rect 218298 183922 220554 183978
rect 220610 183922 220678 183978
rect 220734 183922 220802 183978
rect 220858 183922 220926 183978
rect 220982 183922 248838 183978
rect 248894 183922 248962 183978
rect 249018 183922 251274 183978
rect 251330 183922 251398 183978
rect 251454 183922 251522 183978
rect 251578 183922 251646 183978
rect 251702 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 361130 183978
rect 361186 183922 361254 183978
rect 361310 183922 361378 183978
rect 361434 183922 361502 183978
rect 361558 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 404874 183978
rect 404930 183922 404998 183978
rect 405054 183922 405122 183978
rect 405178 183922 405246 183978
rect 405302 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 445812 183978
rect 445868 183922 445936 183978
rect 445992 183922 446060 183978
rect 446116 183922 446184 183978
rect 446240 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 472732 183978
rect 472788 183922 472856 183978
rect 472912 183922 472980 183978
rect 473036 183922 473104 183978
rect 473160 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 557414 183978
rect 557470 183922 557538 183978
rect 557594 183922 557662 183978
rect 557718 183922 557786 183978
rect 557842 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect 185596 175618 218500 175634
rect 185596 175562 185612 175618
rect 185668 175562 218428 175618
rect 218484 175562 218500 175618
rect 185596 175546 218500 175562
rect 188956 173998 221860 174014
rect 188956 173942 188972 173998
rect 189028 173942 221788 173998
rect 221844 173942 221860 173998
rect 188956 173926 221860 173942
rect 160396 173818 203380 173834
rect 160396 173762 160412 173818
rect 160468 173762 203308 173818
rect 203364 173762 203380 173818
rect 160396 173746 203380 173762
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 70674 172350
rect 70730 172294 70798 172350
rect 70854 172294 70922 172350
rect 70978 172294 71046 172350
rect 71102 172294 79878 172350
rect 79934 172294 80002 172350
rect 80058 172294 101394 172350
rect 101450 172294 101518 172350
rect 101574 172294 101642 172350
rect 101698 172294 101766 172350
rect 101822 172294 110598 172350
rect 110654 172294 110722 172350
rect 110778 172294 132114 172350
rect 132170 172294 132238 172350
rect 132294 172294 132362 172350
rect 132418 172294 132486 172350
rect 132542 172294 141318 172350
rect 141374 172294 141442 172350
rect 141498 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 172038 172350
rect 172094 172294 172162 172350
rect 172218 172294 193554 172350
rect 193610 172294 193678 172350
rect 193734 172294 193802 172350
rect 193858 172294 193926 172350
rect 193982 172294 202758 172350
rect 202814 172294 202882 172350
rect 202938 172294 224274 172350
rect 224330 172294 224398 172350
rect 224454 172294 224522 172350
rect 224578 172294 224646 172350
rect 224702 172294 233478 172350
rect 233534 172294 233602 172350
rect 233658 172294 254994 172350
rect 255050 172294 255118 172350
rect 255174 172294 255242 172350
rect 255298 172294 255366 172350
rect 255422 172294 264198 172350
rect 264254 172294 264322 172350
rect 264378 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 361930 172350
rect 361986 172294 362054 172350
rect 362110 172294 362178 172350
rect 362234 172294 362302 172350
rect 362358 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 446612 172350
rect 446668 172294 446736 172350
rect 446792 172294 446860 172350
rect 446916 172294 446984 172350
rect 447040 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 471932 172350
rect 471988 172294 472056 172350
rect 472112 172294 472180 172350
rect 472236 172294 472304 172350
rect 472360 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 556614 172350
rect 556670 172294 556738 172350
rect 556794 172294 556862 172350
rect 556918 172294 556986 172350
rect 557042 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 70674 172226
rect 70730 172170 70798 172226
rect 70854 172170 70922 172226
rect 70978 172170 71046 172226
rect 71102 172170 79878 172226
rect 79934 172170 80002 172226
rect 80058 172170 101394 172226
rect 101450 172170 101518 172226
rect 101574 172170 101642 172226
rect 101698 172170 101766 172226
rect 101822 172170 110598 172226
rect 110654 172170 110722 172226
rect 110778 172170 132114 172226
rect 132170 172170 132238 172226
rect 132294 172170 132362 172226
rect 132418 172170 132486 172226
rect 132542 172170 141318 172226
rect 141374 172170 141442 172226
rect 141498 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 172038 172226
rect 172094 172170 172162 172226
rect 172218 172170 193554 172226
rect 193610 172170 193678 172226
rect 193734 172170 193802 172226
rect 193858 172170 193926 172226
rect 193982 172170 202758 172226
rect 202814 172170 202882 172226
rect 202938 172170 224274 172226
rect 224330 172170 224398 172226
rect 224454 172170 224522 172226
rect 224578 172170 224646 172226
rect 224702 172170 233478 172226
rect 233534 172170 233602 172226
rect 233658 172170 254994 172226
rect 255050 172170 255118 172226
rect 255174 172170 255242 172226
rect 255298 172170 255366 172226
rect 255422 172170 264198 172226
rect 264254 172170 264322 172226
rect 264378 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 361930 172226
rect 361986 172170 362054 172226
rect 362110 172170 362178 172226
rect 362234 172170 362302 172226
rect 362358 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 446612 172226
rect 446668 172170 446736 172226
rect 446792 172170 446860 172226
rect 446916 172170 446984 172226
rect 447040 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 471932 172226
rect 471988 172170 472056 172226
rect 472112 172170 472180 172226
rect 472236 172170 472304 172226
rect 472360 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 556614 172226
rect 556670 172170 556738 172226
rect 556794 172170 556862 172226
rect 556918 172170 556986 172226
rect 557042 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 70674 172102
rect 70730 172046 70798 172102
rect 70854 172046 70922 172102
rect 70978 172046 71046 172102
rect 71102 172046 79878 172102
rect 79934 172046 80002 172102
rect 80058 172046 101394 172102
rect 101450 172046 101518 172102
rect 101574 172046 101642 172102
rect 101698 172046 101766 172102
rect 101822 172046 110598 172102
rect 110654 172046 110722 172102
rect 110778 172046 132114 172102
rect 132170 172046 132238 172102
rect 132294 172046 132362 172102
rect 132418 172046 132486 172102
rect 132542 172046 141318 172102
rect 141374 172046 141442 172102
rect 141498 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 172038 172102
rect 172094 172046 172162 172102
rect 172218 172046 193554 172102
rect 193610 172046 193678 172102
rect 193734 172046 193802 172102
rect 193858 172046 193926 172102
rect 193982 172046 202758 172102
rect 202814 172046 202882 172102
rect 202938 172046 224274 172102
rect 224330 172046 224398 172102
rect 224454 172046 224522 172102
rect 224578 172046 224646 172102
rect 224702 172046 233478 172102
rect 233534 172046 233602 172102
rect 233658 172046 254994 172102
rect 255050 172046 255118 172102
rect 255174 172046 255242 172102
rect 255298 172046 255366 172102
rect 255422 172046 264198 172102
rect 264254 172046 264322 172102
rect 264378 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 361930 172102
rect 361986 172046 362054 172102
rect 362110 172046 362178 172102
rect 362234 172046 362302 172102
rect 362358 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 446612 172102
rect 446668 172046 446736 172102
rect 446792 172046 446860 172102
rect 446916 172046 446984 172102
rect 447040 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 471932 172102
rect 471988 172046 472056 172102
rect 472112 172046 472180 172102
rect 472236 172046 472304 172102
rect 472360 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 556614 172102
rect 556670 172046 556738 172102
rect 556794 172046 556862 172102
rect 556918 172046 556986 172102
rect 557042 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 70674 171978
rect 70730 171922 70798 171978
rect 70854 171922 70922 171978
rect 70978 171922 71046 171978
rect 71102 171922 79878 171978
rect 79934 171922 80002 171978
rect 80058 171922 101394 171978
rect 101450 171922 101518 171978
rect 101574 171922 101642 171978
rect 101698 171922 101766 171978
rect 101822 171922 110598 171978
rect 110654 171922 110722 171978
rect 110778 171922 132114 171978
rect 132170 171922 132238 171978
rect 132294 171922 132362 171978
rect 132418 171922 132486 171978
rect 132542 171922 141318 171978
rect 141374 171922 141442 171978
rect 141498 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 172038 171978
rect 172094 171922 172162 171978
rect 172218 171922 193554 171978
rect 193610 171922 193678 171978
rect 193734 171922 193802 171978
rect 193858 171922 193926 171978
rect 193982 171922 202758 171978
rect 202814 171922 202882 171978
rect 202938 171922 224274 171978
rect 224330 171922 224398 171978
rect 224454 171922 224522 171978
rect 224578 171922 224646 171978
rect 224702 171922 233478 171978
rect 233534 171922 233602 171978
rect 233658 171922 254994 171978
rect 255050 171922 255118 171978
rect 255174 171922 255242 171978
rect 255298 171922 255366 171978
rect 255422 171922 264198 171978
rect 264254 171922 264322 171978
rect 264378 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 361930 171978
rect 361986 171922 362054 171978
rect 362110 171922 362178 171978
rect 362234 171922 362302 171978
rect 362358 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 446612 171978
rect 446668 171922 446736 171978
rect 446792 171922 446860 171978
rect 446916 171922 446984 171978
rect 447040 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 471932 171978
rect 471988 171922 472056 171978
rect 472112 171922 472180 171978
rect 472236 171922 472304 171978
rect 472360 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 556614 171978
rect 556670 171922 556738 171978
rect 556794 171922 556862 171978
rect 556918 171922 556986 171978
rect 557042 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect 192316 170758 215140 170774
rect 192316 170702 192332 170758
rect 192388 170702 215068 170758
rect 215124 170702 215140 170758
rect 192316 170686 215140 170702
rect 167900 170578 200804 170594
rect 167900 170522 167916 170578
rect 167972 170522 200732 170578
rect 200788 170522 200804 170578
rect 167900 170506 200804 170522
rect 195676 168958 213460 168974
rect 195676 168902 195692 168958
rect 195748 168902 213388 168958
rect 213444 168902 213460 168958
rect 195676 168886 213460 168902
rect 157036 168778 208420 168794
rect 157036 168722 157052 168778
rect 157108 168722 208348 168778
rect 208404 168722 208420 168778
rect 157036 168706 208420 168722
rect 152108 167338 198340 167354
rect 152108 167282 152124 167338
rect 152180 167282 198268 167338
rect 198324 167282 198340 167338
rect 152108 167266 198340 167282
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 64518 166350
rect 64574 166294 64642 166350
rect 64698 166294 66954 166350
rect 67010 166294 67078 166350
rect 67134 166294 67202 166350
rect 67258 166294 67326 166350
rect 67382 166294 95238 166350
rect 95294 166294 95362 166350
rect 95418 166294 97674 166350
rect 97730 166294 97798 166350
rect 97854 166294 97922 166350
rect 97978 166294 98046 166350
rect 98102 166294 125958 166350
rect 126014 166294 126082 166350
rect 126138 166294 128394 166350
rect 128450 166294 128518 166350
rect 128574 166294 128642 166350
rect 128698 166294 128766 166350
rect 128822 166294 156678 166350
rect 156734 166294 156802 166350
rect 156858 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 187398 166350
rect 187454 166294 187522 166350
rect 187578 166294 189834 166350
rect 189890 166294 189958 166350
rect 190014 166294 190082 166350
rect 190138 166294 190206 166350
rect 190262 166294 218118 166350
rect 218174 166294 218242 166350
rect 218298 166294 248838 166350
rect 248894 166294 248962 166350
rect 249018 166294 251274 166350
rect 251330 166294 251398 166350
rect 251454 166294 251522 166350
rect 251578 166294 251646 166350
rect 251702 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 361130 166350
rect 361186 166294 361254 166350
rect 361310 166294 361378 166350
rect 361434 166294 361502 166350
rect 361558 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 445812 166350
rect 445868 166294 445936 166350
rect 445992 166294 446060 166350
rect 446116 166294 446184 166350
rect 446240 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 472732 166350
rect 472788 166294 472856 166350
rect 472912 166294 472980 166350
rect 473036 166294 473104 166350
rect 473160 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 557414 166350
rect 557470 166294 557538 166350
rect 557594 166294 557662 166350
rect 557718 166294 557786 166350
rect 557842 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 64518 166226
rect 64574 166170 64642 166226
rect 64698 166170 66954 166226
rect 67010 166170 67078 166226
rect 67134 166170 67202 166226
rect 67258 166170 67326 166226
rect 67382 166170 95238 166226
rect 95294 166170 95362 166226
rect 95418 166170 97674 166226
rect 97730 166170 97798 166226
rect 97854 166170 97922 166226
rect 97978 166170 98046 166226
rect 98102 166170 125958 166226
rect 126014 166170 126082 166226
rect 126138 166170 128394 166226
rect 128450 166170 128518 166226
rect 128574 166170 128642 166226
rect 128698 166170 128766 166226
rect 128822 166170 156678 166226
rect 156734 166170 156802 166226
rect 156858 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 187398 166226
rect 187454 166170 187522 166226
rect 187578 166170 189834 166226
rect 189890 166170 189958 166226
rect 190014 166170 190082 166226
rect 190138 166170 190206 166226
rect 190262 166170 218118 166226
rect 218174 166170 218242 166226
rect 218298 166170 248838 166226
rect 248894 166170 248962 166226
rect 249018 166170 251274 166226
rect 251330 166170 251398 166226
rect 251454 166170 251522 166226
rect 251578 166170 251646 166226
rect 251702 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 361130 166226
rect 361186 166170 361254 166226
rect 361310 166170 361378 166226
rect 361434 166170 361502 166226
rect 361558 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 445812 166226
rect 445868 166170 445936 166226
rect 445992 166170 446060 166226
rect 446116 166170 446184 166226
rect 446240 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 472732 166226
rect 472788 166170 472856 166226
rect 472912 166170 472980 166226
rect 473036 166170 473104 166226
rect 473160 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 557414 166226
rect 557470 166170 557538 166226
rect 557594 166170 557662 166226
rect 557718 166170 557786 166226
rect 557842 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 64518 166102
rect 64574 166046 64642 166102
rect 64698 166046 66954 166102
rect 67010 166046 67078 166102
rect 67134 166046 67202 166102
rect 67258 166046 67326 166102
rect 67382 166046 95238 166102
rect 95294 166046 95362 166102
rect 95418 166046 97674 166102
rect 97730 166046 97798 166102
rect 97854 166046 97922 166102
rect 97978 166046 98046 166102
rect 98102 166046 125958 166102
rect 126014 166046 126082 166102
rect 126138 166046 128394 166102
rect 128450 166046 128518 166102
rect 128574 166046 128642 166102
rect 128698 166046 128766 166102
rect 128822 166046 156678 166102
rect 156734 166046 156802 166102
rect 156858 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 187398 166102
rect 187454 166046 187522 166102
rect 187578 166046 189834 166102
rect 189890 166046 189958 166102
rect 190014 166046 190082 166102
rect 190138 166046 190206 166102
rect 190262 166046 218118 166102
rect 218174 166046 218242 166102
rect 218298 166046 248838 166102
rect 248894 166046 248962 166102
rect 249018 166046 251274 166102
rect 251330 166046 251398 166102
rect 251454 166046 251522 166102
rect 251578 166046 251646 166102
rect 251702 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 361130 166102
rect 361186 166046 361254 166102
rect 361310 166046 361378 166102
rect 361434 166046 361502 166102
rect 361558 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 445812 166102
rect 445868 166046 445936 166102
rect 445992 166046 446060 166102
rect 446116 166046 446184 166102
rect 446240 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 472732 166102
rect 472788 166046 472856 166102
rect 472912 166046 472980 166102
rect 473036 166046 473104 166102
rect 473160 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 557414 166102
rect 557470 166046 557538 166102
rect 557594 166046 557662 166102
rect 557718 166046 557786 166102
rect 557842 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 64518 165978
rect 64574 165922 64642 165978
rect 64698 165922 66954 165978
rect 67010 165922 67078 165978
rect 67134 165922 67202 165978
rect 67258 165922 67326 165978
rect 67382 165922 95238 165978
rect 95294 165922 95362 165978
rect 95418 165922 97674 165978
rect 97730 165922 97798 165978
rect 97854 165922 97922 165978
rect 97978 165922 98046 165978
rect 98102 165922 125958 165978
rect 126014 165922 126082 165978
rect 126138 165922 128394 165978
rect 128450 165922 128518 165978
rect 128574 165922 128642 165978
rect 128698 165922 128766 165978
rect 128822 165922 156678 165978
rect 156734 165922 156802 165978
rect 156858 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 187398 165978
rect 187454 165922 187522 165978
rect 187578 165922 189834 165978
rect 189890 165922 189958 165978
rect 190014 165922 190082 165978
rect 190138 165922 190206 165978
rect 190262 165922 218118 165978
rect 218174 165922 218242 165978
rect 218298 165922 248838 165978
rect 248894 165922 248962 165978
rect 249018 165922 251274 165978
rect 251330 165922 251398 165978
rect 251454 165922 251522 165978
rect 251578 165922 251646 165978
rect 251702 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 361130 165978
rect 361186 165922 361254 165978
rect 361310 165922 361378 165978
rect 361434 165922 361502 165978
rect 361558 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 445812 165978
rect 445868 165922 445936 165978
rect 445992 165922 446060 165978
rect 446116 165922 446184 165978
rect 446240 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 472732 165978
rect 472788 165922 472856 165978
rect 472912 165922 472980 165978
rect 473036 165922 473104 165978
rect 473160 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 557414 165978
rect 557470 165922 557538 165978
rect 557594 165922 557662 165978
rect 557718 165922 557786 165978
rect 557842 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 70674 154350
rect 70730 154294 70798 154350
rect 70854 154294 70922 154350
rect 70978 154294 71046 154350
rect 71102 154294 101394 154350
rect 101450 154294 101518 154350
rect 101574 154294 101642 154350
rect 101698 154294 101766 154350
rect 101822 154294 132114 154350
rect 132170 154294 132238 154350
rect 132294 154294 132362 154350
rect 132418 154294 132486 154350
rect 132542 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 193554 154350
rect 193610 154294 193678 154350
rect 193734 154294 193802 154350
rect 193858 154294 193926 154350
rect 193982 154294 224274 154350
rect 224330 154294 224398 154350
rect 224454 154294 224522 154350
rect 224578 154294 224646 154350
rect 224702 154294 254994 154350
rect 255050 154294 255118 154350
rect 255174 154294 255242 154350
rect 255298 154294 255366 154350
rect 255422 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 70674 154226
rect 70730 154170 70798 154226
rect 70854 154170 70922 154226
rect 70978 154170 71046 154226
rect 71102 154170 101394 154226
rect 101450 154170 101518 154226
rect 101574 154170 101642 154226
rect 101698 154170 101766 154226
rect 101822 154170 132114 154226
rect 132170 154170 132238 154226
rect 132294 154170 132362 154226
rect 132418 154170 132486 154226
rect 132542 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 193554 154226
rect 193610 154170 193678 154226
rect 193734 154170 193802 154226
rect 193858 154170 193926 154226
rect 193982 154170 224274 154226
rect 224330 154170 224398 154226
rect 224454 154170 224522 154226
rect 224578 154170 224646 154226
rect 224702 154170 254994 154226
rect 255050 154170 255118 154226
rect 255174 154170 255242 154226
rect 255298 154170 255366 154226
rect 255422 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 70674 154102
rect 70730 154046 70798 154102
rect 70854 154046 70922 154102
rect 70978 154046 71046 154102
rect 71102 154046 101394 154102
rect 101450 154046 101518 154102
rect 101574 154046 101642 154102
rect 101698 154046 101766 154102
rect 101822 154046 132114 154102
rect 132170 154046 132238 154102
rect 132294 154046 132362 154102
rect 132418 154046 132486 154102
rect 132542 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 193554 154102
rect 193610 154046 193678 154102
rect 193734 154046 193802 154102
rect 193858 154046 193926 154102
rect 193982 154046 224274 154102
rect 224330 154046 224398 154102
rect 224454 154046 224522 154102
rect 224578 154046 224646 154102
rect 224702 154046 254994 154102
rect 255050 154046 255118 154102
rect 255174 154046 255242 154102
rect 255298 154046 255366 154102
rect 255422 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 70674 153978
rect 70730 153922 70798 153978
rect 70854 153922 70922 153978
rect 70978 153922 71046 153978
rect 71102 153922 101394 153978
rect 101450 153922 101518 153978
rect 101574 153922 101642 153978
rect 101698 153922 101766 153978
rect 101822 153922 132114 153978
rect 132170 153922 132238 153978
rect 132294 153922 132362 153978
rect 132418 153922 132486 153978
rect 132542 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 193554 153978
rect 193610 153922 193678 153978
rect 193734 153922 193802 153978
rect 193858 153922 193926 153978
rect 193982 153922 224274 153978
rect 224330 153922 224398 153978
rect 224454 153922 224522 153978
rect 224578 153922 224646 153978
rect 224702 153922 254994 153978
rect 255050 153922 255118 153978
rect 255174 153922 255242 153978
rect 255298 153922 255366 153978
rect 255422 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 66954 148350
rect 67010 148294 67078 148350
rect 67134 148294 67202 148350
rect 67258 148294 67326 148350
rect 67382 148294 97674 148350
rect 97730 148294 97798 148350
rect 97854 148294 97922 148350
rect 97978 148294 98046 148350
rect 98102 148294 128394 148350
rect 128450 148294 128518 148350
rect 128574 148294 128642 148350
rect 128698 148294 128766 148350
rect 128822 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 189834 148350
rect 189890 148294 189958 148350
rect 190014 148294 190082 148350
rect 190138 148294 190206 148350
rect 190262 148294 220554 148350
rect 220610 148294 220678 148350
rect 220734 148294 220802 148350
rect 220858 148294 220926 148350
rect 220982 148294 251274 148350
rect 251330 148294 251398 148350
rect 251454 148294 251522 148350
rect 251578 148294 251646 148350
rect 251702 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 466314 148350
rect 466370 148294 466438 148350
rect 466494 148294 466562 148350
rect 466618 148294 466686 148350
rect 466742 148294 497034 148350
rect 497090 148294 497158 148350
rect 497214 148294 497282 148350
rect 497338 148294 497406 148350
rect 497462 148294 527754 148350
rect 527810 148294 527878 148350
rect 527934 148294 528002 148350
rect 528058 148294 528126 148350
rect 528182 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 66954 148226
rect 67010 148170 67078 148226
rect 67134 148170 67202 148226
rect 67258 148170 67326 148226
rect 67382 148170 97674 148226
rect 97730 148170 97798 148226
rect 97854 148170 97922 148226
rect 97978 148170 98046 148226
rect 98102 148170 128394 148226
rect 128450 148170 128518 148226
rect 128574 148170 128642 148226
rect 128698 148170 128766 148226
rect 128822 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 189834 148226
rect 189890 148170 189958 148226
rect 190014 148170 190082 148226
rect 190138 148170 190206 148226
rect 190262 148170 220554 148226
rect 220610 148170 220678 148226
rect 220734 148170 220802 148226
rect 220858 148170 220926 148226
rect 220982 148170 251274 148226
rect 251330 148170 251398 148226
rect 251454 148170 251522 148226
rect 251578 148170 251646 148226
rect 251702 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 466314 148226
rect 466370 148170 466438 148226
rect 466494 148170 466562 148226
rect 466618 148170 466686 148226
rect 466742 148170 497034 148226
rect 497090 148170 497158 148226
rect 497214 148170 497282 148226
rect 497338 148170 497406 148226
rect 497462 148170 527754 148226
rect 527810 148170 527878 148226
rect 527934 148170 528002 148226
rect 528058 148170 528126 148226
rect 528182 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 66954 148102
rect 67010 148046 67078 148102
rect 67134 148046 67202 148102
rect 67258 148046 67326 148102
rect 67382 148046 97674 148102
rect 97730 148046 97798 148102
rect 97854 148046 97922 148102
rect 97978 148046 98046 148102
rect 98102 148046 128394 148102
rect 128450 148046 128518 148102
rect 128574 148046 128642 148102
rect 128698 148046 128766 148102
rect 128822 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 189834 148102
rect 189890 148046 189958 148102
rect 190014 148046 190082 148102
rect 190138 148046 190206 148102
rect 190262 148046 220554 148102
rect 220610 148046 220678 148102
rect 220734 148046 220802 148102
rect 220858 148046 220926 148102
rect 220982 148046 251274 148102
rect 251330 148046 251398 148102
rect 251454 148046 251522 148102
rect 251578 148046 251646 148102
rect 251702 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 466314 148102
rect 466370 148046 466438 148102
rect 466494 148046 466562 148102
rect 466618 148046 466686 148102
rect 466742 148046 497034 148102
rect 497090 148046 497158 148102
rect 497214 148046 497282 148102
rect 497338 148046 497406 148102
rect 497462 148046 527754 148102
rect 527810 148046 527878 148102
rect 527934 148046 528002 148102
rect 528058 148046 528126 148102
rect 528182 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 66954 147978
rect 67010 147922 67078 147978
rect 67134 147922 67202 147978
rect 67258 147922 67326 147978
rect 67382 147922 97674 147978
rect 97730 147922 97798 147978
rect 97854 147922 97922 147978
rect 97978 147922 98046 147978
rect 98102 147922 128394 147978
rect 128450 147922 128518 147978
rect 128574 147922 128642 147978
rect 128698 147922 128766 147978
rect 128822 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 189834 147978
rect 189890 147922 189958 147978
rect 190014 147922 190082 147978
rect 190138 147922 190206 147978
rect 190262 147922 220554 147978
rect 220610 147922 220678 147978
rect 220734 147922 220802 147978
rect 220858 147922 220926 147978
rect 220982 147922 251274 147978
rect 251330 147922 251398 147978
rect 251454 147922 251522 147978
rect 251578 147922 251646 147978
rect 251702 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 466314 147978
rect 466370 147922 466438 147978
rect 466494 147922 466562 147978
rect 466618 147922 466686 147978
rect 466742 147922 497034 147978
rect 497090 147922 497158 147978
rect 497214 147922 497282 147978
rect 497338 147922 497406 147978
rect 497462 147922 527754 147978
rect 527810 147922 527878 147978
rect 527934 147922 528002 147978
rect 528058 147922 528126 147978
rect 528182 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect 62172 142678 119380 142694
rect 62172 142622 62188 142678
rect 62244 142622 62748 142678
rect 62804 142622 119308 142678
rect 119364 142622 119380 142678
rect 62172 142606 119380 142622
rect 144716 142678 243644 142694
rect 144716 142622 144732 142678
rect 144788 142622 243644 142678
rect 144716 142606 243644 142622
rect 418332 142678 499060 142694
rect 418332 142622 418348 142678
rect 418404 142622 498988 142678
rect 499044 142622 499060 142678
rect 418332 142606 499060 142622
rect 63740 142318 131028 142334
rect 63740 142262 63756 142318
rect 63812 142262 130956 142318
rect 131012 142262 131028 142318
rect 63740 142246 131028 142262
rect 243556 142154 243644 142606
rect 349396 142498 544756 142514
rect 349396 142442 444668 142498
rect 444724 142442 474572 142498
rect 474628 142442 544684 142498
rect 544740 142442 544756 142498
rect 349396 142426 544756 142442
rect 349396 142154 349484 142426
rect 445548 142318 472068 142334
rect 445548 142262 445564 142318
rect 445620 142262 471996 142318
rect 472052 142262 472068 142318
rect 445548 142246 472068 142262
rect 84908 142138 164516 142154
rect 84908 142082 84924 142138
rect 84980 142082 164444 142138
rect 164500 142082 164516 142138
rect 84908 142066 164516 142082
rect 243556 142138 349484 142154
rect 243556 142082 244636 142138
rect 244692 142082 304780 142138
rect 304836 142082 344652 142138
rect 344708 142082 349484 142138
rect 243556 142066 349484 142082
rect 119292 141958 418420 141974
rect 119292 141902 119308 141958
rect 119364 141902 219324 141958
rect 219380 141902 319228 141958
rect 319284 141902 330876 141958
rect 330932 141902 418348 141958
rect 418404 141902 418420 141958
rect 119292 141886 418420 141902
rect 484412 141958 534676 141974
rect 484412 141902 484428 141958
rect 484484 141902 534604 141958
rect 534660 141902 534676 141958
rect 484412 141886 534676 141902
rect 114700 141058 505668 141074
rect 114700 141002 114716 141058
rect 114772 141002 214620 141058
rect 214676 141002 314636 141058
rect 314692 141002 333452 141058
rect 333508 141002 414652 141058
rect 414708 141002 505596 141058
rect 505652 141002 505668 141058
rect 114700 140986 505668 141002
rect 145388 140878 245492 140894
rect 145388 140822 145404 140878
rect 145460 140822 245420 140878
rect 245476 140822 245492 140878
rect 145388 140806 245492 140822
rect 303980 140878 341028 140894
rect 303980 140822 303996 140878
rect 304052 140822 340956 140878
rect 341012 140822 341028 140878
rect 303980 140806 341028 140822
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 70674 136350
rect 70730 136294 70798 136350
rect 70854 136294 70922 136350
rect 70978 136294 71046 136350
rect 71102 136294 101394 136350
rect 101450 136294 101518 136350
rect 101574 136294 101642 136350
rect 101698 136294 101766 136350
rect 101822 136294 132114 136350
rect 132170 136294 132238 136350
rect 132294 136294 132362 136350
rect 132418 136294 132486 136350
rect 132542 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 193554 136350
rect 193610 136294 193678 136350
rect 193734 136294 193802 136350
rect 193858 136294 193926 136350
rect 193982 136294 224274 136350
rect 224330 136294 224398 136350
rect 224454 136294 224522 136350
rect 224578 136294 224646 136350
rect 224702 136294 254994 136350
rect 255050 136294 255118 136350
rect 255174 136294 255242 136350
rect 255298 136294 255366 136350
rect 255422 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 470034 136350
rect 470090 136294 470158 136350
rect 470214 136294 470282 136350
rect 470338 136294 470406 136350
rect 470462 136294 500754 136350
rect 500810 136294 500878 136350
rect 500934 136294 501002 136350
rect 501058 136294 501126 136350
rect 501182 136294 531474 136350
rect 531530 136294 531598 136350
rect 531654 136294 531722 136350
rect 531778 136294 531846 136350
rect 531902 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 70674 136226
rect 70730 136170 70798 136226
rect 70854 136170 70922 136226
rect 70978 136170 71046 136226
rect 71102 136170 101394 136226
rect 101450 136170 101518 136226
rect 101574 136170 101642 136226
rect 101698 136170 101766 136226
rect 101822 136170 132114 136226
rect 132170 136170 132238 136226
rect 132294 136170 132362 136226
rect 132418 136170 132486 136226
rect 132542 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 193554 136226
rect 193610 136170 193678 136226
rect 193734 136170 193802 136226
rect 193858 136170 193926 136226
rect 193982 136170 224274 136226
rect 224330 136170 224398 136226
rect 224454 136170 224522 136226
rect 224578 136170 224646 136226
rect 224702 136170 254994 136226
rect 255050 136170 255118 136226
rect 255174 136170 255242 136226
rect 255298 136170 255366 136226
rect 255422 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 470034 136226
rect 470090 136170 470158 136226
rect 470214 136170 470282 136226
rect 470338 136170 470406 136226
rect 470462 136170 500754 136226
rect 500810 136170 500878 136226
rect 500934 136170 501002 136226
rect 501058 136170 501126 136226
rect 501182 136170 531474 136226
rect 531530 136170 531598 136226
rect 531654 136170 531722 136226
rect 531778 136170 531846 136226
rect 531902 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 70674 136102
rect 70730 136046 70798 136102
rect 70854 136046 70922 136102
rect 70978 136046 71046 136102
rect 71102 136046 101394 136102
rect 101450 136046 101518 136102
rect 101574 136046 101642 136102
rect 101698 136046 101766 136102
rect 101822 136046 132114 136102
rect 132170 136046 132238 136102
rect 132294 136046 132362 136102
rect 132418 136046 132486 136102
rect 132542 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 193554 136102
rect 193610 136046 193678 136102
rect 193734 136046 193802 136102
rect 193858 136046 193926 136102
rect 193982 136046 224274 136102
rect 224330 136046 224398 136102
rect 224454 136046 224522 136102
rect 224578 136046 224646 136102
rect 224702 136046 254994 136102
rect 255050 136046 255118 136102
rect 255174 136046 255242 136102
rect 255298 136046 255366 136102
rect 255422 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 470034 136102
rect 470090 136046 470158 136102
rect 470214 136046 470282 136102
rect 470338 136046 470406 136102
rect 470462 136046 500754 136102
rect 500810 136046 500878 136102
rect 500934 136046 501002 136102
rect 501058 136046 501126 136102
rect 501182 136046 531474 136102
rect 531530 136046 531598 136102
rect 531654 136046 531722 136102
rect 531778 136046 531846 136102
rect 531902 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 70674 135978
rect 70730 135922 70798 135978
rect 70854 135922 70922 135978
rect 70978 135922 71046 135978
rect 71102 135922 101394 135978
rect 101450 135922 101518 135978
rect 101574 135922 101642 135978
rect 101698 135922 101766 135978
rect 101822 135922 132114 135978
rect 132170 135922 132238 135978
rect 132294 135922 132362 135978
rect 132418 135922 132486 135978
rect 132542 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 193554 135978
rect 193610 135922 193678 135978
rect 193734 135922 193802 135978
rect 193858 135922 193926 135978
rect 193982 135922 224274 135978
rect 224330 135922 224398 135978
rect 224454 135922 224522 135978
rect 224578 135922 224646 135978
rect 224702 135922 254994 135978
rect 255050 135922 255118 135978
rect 255174 135922 255242 135978
rect 255298 135922 255366 135978
rect 255422 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 470034 135978
rect 470090 135922 470158 135978
rect 470214 135922 470282 135978
rect 470338 135922 470406 135978
rect 470462 135922 500754 135978
rect 500810 135922 500878 135978
rect 500934 135922 501002 135978
rect 501058 135922 501126 135978
rect 501182 135922 531474 135978
rect 531530 135922 531598 135978
rect 531654 135922 531722 135978
rect 531778 135922 531846 135978
rect 531902 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 61130 130350
rect 61186 130294 61254 130350
rect 61310 130294 61378 130350
rect 61434 130294 61502 130350
rect 61558 130294 66954 130350
rect 67010 130294 67078 130350
rect 67134 130294 67202 130350
rect 67258 130294 67326 130350
rect 67382 130294 97674 130350
rect 97730 130294 97798 130350
rect 97854 130294 97922 130350
rect 97978 130294 98046 130350
rect 98102 130294 128394 130350
rect 128450 130294 128518 130350
rect 128574 130294 128642 130350
rect 128698 130294 128766 130350
rect 128822 130294 145812 130350
rect 145868 130294 145936 130350
rect 145992 130294 146060 130350
rect 146116 130294 146184 130350
rect 146240 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 161130 130350
rect 161186 130294 161254 130350
rect 161310 130294 161378 130350
rect 161434 130294 161502 130350
rect 161558 130294 189834 130350
rect 189890 130294 189958 130350
rect 190014 130294 190082 130350
rect 190138 130294 190206 130350
rect 190262 130294 220554 130350
rect 220610 130294 220678 130350
rect 220734 130294 220802 130350
rect 220858 130294 220926 130350
rect 220982 130294 245812 130350
rect 245868 130294 245936 130350
rect 245992 130294 246060 130350
rect 246116 130294 246184 130350
rect 246240 130294 251274 130350
rect 251330 130294 251398 130350
rect 251454 130294 251522 130350
rect 251578 130294 251646 130350
rect 251702 130294 261130 130350
rect 261186 130294 261254 130350
rect 261310 130294 261378 130350
rect 261434 130294 261502 130350
rect 261558 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 345812 130350
rect 345868 130294 345936 130350
rect 345992 130294 346060 130350
rect 346116 130294 346184 130350
rect 346240 130294 361130 130350
rect 361186 130294 361254 130350
rect 361310 130294 361378 130350
rect 361434 130294 361502 130350
rect 361558 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 445812 130350
rect 445868 130294 445936 130350
rect 445992 130294 446060 130350
rect 446116 130294 446184 130350
rect 446240 130294 461130 130350
rect 461186 130294 461254 130350
rect 461310 130294 461378 130350
rect 461434 130294 461502 130350
rect 461558 130294 466314 130350
rect 466370 130294 466438 130350
rect 466494 130294 466562 130350
rect 466618 130294 466686 130350
rect 466742 130294 497034 130350
rect 497090 130294 497158 130350
rect 497214 130294 497282 130350
rect 497338 130294 497406 130350
rect 497462 130294 527754 130350
rect 527810 130294 527878 130350
rect 527934 130294 528002 130350
rect 528058 130294 528126 130350
rect 528182 130294 545812 130350
rect 545868 130294 545936 130350
rect 545992 130294 546060 130350
rect 546116 130294 546184 130350
rect 546240 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 61130 130226
rect 61186 130170 61254 130226
rect 61310 130170 61378 130226
rect 61434 130170 61502 130226
rect 61558 130170 66954 130226
rect 67010 130170 67078 130226
rect 67134 130170 67202 130226
rect 67258 130170 67326 130226
rect 67382 130170 97674 130226
rect 97730 130170 97798 130226
rect 97854 130170 97922 130226
rect 97978 130170 98046 130226
rect 98102 130170 128394 130226
rect 128450 130170 128518 130226
rect 128574 130170 128642 130226
rect 128698 130170 128766 130226
rect 128822 130170 145812 130226
rect 145868 130170 145936 130226
rect 145992 130170 146060 130226
rect 146116 130170 146184 130226
rect 146240 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 161130 130226
rect 161186 130170 161254 130226
rect 161310 130170 161378 130226
rect 161434 130170 161502 130226
rect 161558 130170 189834 130226
rect 189890 130170 189958 130226
rect 190014 130170 190082 130226
rect 190138 130170 190206 130226
rect 190262 130170 220554 130226
rect 220610 130170 220678 130226
rect 220734 130170 220802 130226
rect 220858 130170 220926 130226
rect 220982 130170 245812 130226
rect 245868 130170 245936 130226
rect 245992 130170 246060 130226
rect 246116 130170 246184 130226
rect 246240 130170 251274 130226
rect 251330 130170 251398 130226
rect 251454 130170 251522 130226
rect 251578 130170 251646 130226
rect 251702 130170 261130 130226
rect 261186 130170 261254 130226
rect 261310 130170 261378 130226
rect 261434 130170 261502 130226
rect 261558 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 345812 130226
rect 345868 130170 345936 130226
rect 345992 130170 346060 130226
rect 346116 130170 346184 130226
rect 346240 130170 361130 130226
rect 361186 130170 361254 130226
rect 361310 130170 361378 130226
rect 361434 130170 361502 130226
rect 361558 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 445812 130226
rect 445868 130170 445936 130226
rect 445992 130170 446060 130226
rect 446116 130170 446184 130226
rect 446240 130170 461130 130226
rect 461186 130170 461254 130226
rect 461310 130170 461378 130226
rect 461434 130170 461502 130226
rect 461558 130170 466314 130226
rect 466370 130170 466438 130226
rect 466494 130170 466562 130226
rect 466618 130170 466686 130226
rect 466742 130170 497034 130226
rect 497090 130170 497158 130226
rect 497214 130170 497282 130226
rect 497338 130170 497406 130226
rect 497462 130170 527754 130226
rect 527810 130170 527878 130226
rect 527934 130170 528002 130226
rect 528058 130170 528126 130226
rect 528182 130170 545812 130226
rect 545868 130170 545936 130226
rect 545992 130170 546060 130226
rect 546116 130170 546184 130226
rect 546240 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 61130 130102
rect 61186 130046 61254 130102
rect 61310 130046 61378 130102
rect 61434 130046 61502 130102
rect 61558 130046 66954 130102
rect 67010 130046 67078 130102
rect 67134 130046 67202 130102
rect 67258 130046 67326 130102
rect 67382 130046 97674 130102
rect 97730 130046 97798 130102
rect 97854 130046 97922 130102
rect 97978 130046 98046 130102
rect 98102 130046 128394 130102
rect 128450 130046 128518 130102
rect 128574 130046 128642 130102
rect 128698 130046 128766 130102
rect 128822 130046 145812 130102
rect 145868 130046 145936 130102
rect 145992 130046 146060 130102
rect 146116 130046 146184 130102
rect 146240 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 161130 130102
rect 161186 130046 161254 130102
rect 161310 130046 161378 130102
rect 161434 130046 161502 130102
rect 161558 130046 189834 130102
rect 189890 130046 189958 130102
rect 190014 130046 190082 130102
rect 190138 130046 190206 130102
rect 190262 130046 220554 130102
rect 220610 130046 220678 130102
rect 220734 130046 220802 130102
rect 220858 130046 220926 130102
rect 220982 130046 245812 130102
rect 245868 130046 245936 130102
rect 245992 130046 246060 130102
rect 246116 130046 246184 130102
rect 246240 130046 251274 130102
rect 251330 130046 251398 130102
rect 251454 130046 251522 130102
rect 251578 130046 251646 130102
rect 251702 130046 261130 130102
rect 261186 130046 261254 130102
rect 261310 130046 261378 130102
rect 261434 130046 261502 130102
rect 261558 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 345812 130102
rect 345868 130046 345936 130102
rect 345992 130046 346060 130102
rect 346116 130046 346184 130102
rect 346240 130046 361130 130102
rect 361186 130046 361254 130102
rect 361310 130046 361378 130102
rect 361434 130046 361502 130102
rect 361558 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 445812 130102
rect 445868 130046 445936 130102
rect 445992 130046 446060 130102
rect 446116 130046 446184 130102
rect 446240 130046 461130 130102
rect 461186 130046 461254 130102
rect 461310 130046 461378 130102
rect 461434 130046 461502 130102
rect 461558 130046 466314 130102
rect 466370 130046 466438 130102
rect 466494 130046 466562 130102
rect 466618 130046 466686 130102
rect 466742 130046 497034 130102
rect 497090 130046 497158 130102
rect 497214 130046 497282 130102
rect 497338 130046 497406 130102
rect 497462 130046 527754 130102
rect 527810 130046 527878 130102
rect 527934 130046 528002 130102
rect 528058 130046 528126 130102
rect 528182 130046 545812 130102
rect 545868 130046 545936 130102
rect 545992 130046 546060 130102
rect 546116 130046 546184 130102
rect 546240 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 61130 129978
rect 61186 129922 61254 129978
rect 61310 129922 61378 129978
rect 61434 129922 61502 129978
rect 61558 129922 66954 129978
rect 67010 129922 67078 129978
rect 67134 129922 67202 129978
rect 67258 129922 67326 129978
rect 67382 129922 97674 129978
rect 97730 129922 97798 129978
rect 97854 129922 97922 129978
rect 97978 129922 98046 129978
rect 98102 129922 128394 129978
rect 128450 129922 128518 129978
rect 128574 129922 128642 129978
rect 128698 129922 128766 129978
rect 128822 129922 145812 129978
rect 145868 129922 145936 129978
rect 145992 129922 146060 129978
rect 146116 129922 146184 129978
rect 146240 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 161130 129978
rect 161186 129922 161254 129978
rect 161310 129922 161378 129978
rect 161434 129922 161502 129978
rect 161558 129922 189834 129978
rect 189890 129922 189958 129978
rect 190014 129922 190082 129978
rect 190138 129922 190206 129978
rect 190262 129922 220554 129978
rect 220610 129922 220678 129978
rect 220734 129922 220802 129978
rect 220858 129922 220926 129978
rect 220982 129922 245812 129978
rect 245868 129922 245936 129978
rect 245992 129922 246060 129978
rect 246116 129922 246184 129978
rect 246240 129922 251274 129978
rect 251330 129922 251398 129978
rect 251454 129922 251522 129978
rect 251578 129922 251646 129978
rect 251702 129922 261130 129978
rect 261186 129922 261254 129978
rect 261310 129922 261378 129978
rect 261434 129922 261502 129978
rect 261558 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 345812 129978
rect 345868 129922 345936 129978
rect 345992 129922 346060 129978
rect 346116 129922 346184 129978
rect 346240 129922 361130 129978
rect 361186 129922 361254 129978
rect 361310 129922 361378 129978
rect 361434 129922 361502 129978
rect 361558 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 445812 129978
rect 445868 129922 445936 129978
rect 445992 129922 446060 129978
rect 446116 129922 446184 129978
rect 446240 129922 461130 129978
rect 461186 129922 461254 129978
rect 461310 129922 461378 129978
rect 461434 129922 461502 129978
rect 461558 129922 466314 129978
rect 466370 129922 466438 129978
rect 466494 129922 466562 129978
rect 466618 129922 466686 129978
rect 466742 129922 497034 129978
rect 497090 129922 497158 129978
rect 497214 129922 497282 129978
rect 497338 129922 497406 129978
rect 497462 129922 527754 129978
rect 527810 129922 527878 129978
rect 527934 129922 528002 129978
rect 528058 129922 528126 129978
rect 528182 129922 545812 129978
rect 545868 129922 545936 129978
rect 545992 129922 546060 129978
rect 546116 129922 546184 129978
rect 546240 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect 299948 127558 590228 127574
rect 299948 127502 299964 127558
rect 300020 127502 590156 127558
rect 590212 127502 590228 127558
rect 299948 127486 590228 127502
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 61930 118350
rect 61986 118294 62054 118350
rect 62110 118294 62178 118350
rect 62234 118294 62302 118350
rect 62358 118294 70674 118350
rect 70730 118294 70798 118350
rect 70854 118294 70922 118350
rect 70978 118294 71046 118350
rect 71102 118294 101394 118350
rect 101450 118294 101518 118350
rect 101574 118294 101642 118350
rect 101698 118294 101766 118350
rect 101822 118294 132114 118350
rect 132170 118294 132238 118350
rect 132294 118294 132362 118350
rect 132418 118294 132486 118350
rect 132542 118294 146612 118350
rect 146668 118294 146736 118350
rect 146792 118294 146860 118350
rect 146916 118294 146984 118350
rect 147040 118294 161930 118350
rect 161986 118294 162054 118350
rect 162110 118294 162178 118350
rect 162234 118294 162302 118350
rect 162358 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 193554 118350
rect 193610 118294 193678 118350
rect 193734 118294 193802 118350
rect 193858 118294 193926 118350
rect 193982 118294 224274 118350
rect 224330 118294 224398 118350
rect 224454 118294 224522 118350
rect 224578 118294 224646 118350
rect 224702 118294 246612 118350
rect 246668 118294 246736 118350
rect 246792 118294 246860 118350
rect 246916 118294 246984 118350
rect 247040 118294 254994 118350
rect 255050 118294 255118 118350
rect 255174 118294 255242 118350
rect 255298 118294 255366 118350
rect 255422 118294 261930 118350
rect 261986 118294 262054 118350
rect 262110 118294 262178 118350
rect 262234 118294 262302 118350
rect 262358 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 346612 118350
rect 346668 118294 346736 118350
rect 346792 118294 346860 118350
rect 346916 118294 346984 118350
rect 347040 118294 361930 118350
rect 361986 118294 362054 118350
rect 362110 118294 362178 118350
rect 362234 118294 362302 118350
rect 362358 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 446612 118350
rect 446668 118294 446736 118350
rect 446792 118294 446860 118350
rect 446916 118294 446984 118350
rect 447040 118294 461930 118350
rect 461986 118294 462054 118350
rect 462110 118294 462178 118350
rect 462234 118294 462302 118350
rect 462358 118294 470034 118350
rect 470090 118294 470158 118350
rect 470214 118294 470282 118350
rect 470338 118294 470406 118350
rect 470462 118294 500754 118350
rect 500810 118294 500878 118350
rect 500934 118294 501002 118350
rect 501058 118294 501126 118350
rect 501182 118294 531474 118350
rect 531530 118294 531598 118350
rect 531654 118294 531722 118350
rect 531778 118294 531846 118350
rect 531902 118294 546612 118350
rect 546668 118294 546736 118350
rect 546792 118294 546860 118350
rect 546916 118294 546984 118350
rect 547040 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 61930 118226
rect 61986 118170 62054 118226
rect 62110 118170 62178 118226
rect 62234 118170 62302 118226
rect 62358 118170 70674 118226
rect 70730 118170 70798 118226
rect 70854 118170 70922 118226
rect 70978 118170 71046 118226
rect 71102 118170 101394 118226
rect 101450 118170 101518 118226
rect 101574 118170 101642 118226
rect 101698 118170 101766 118226
rect 101822 118170 132114 118226
rect 132170 118170 132238 118226
rect 132294 118170 132362 118226
rect 132418 118170 132486 118226
rect 132542 118170 146612 118226
rect 146668 118170 146736 118226
rect 146792 118170 146860 118226
rect 146916 118170 146984 118226
rect 147040 118170 161930 118226
rect 161986 118170 162054 118226
rect 162110 118170 162178 118226
rect 162234 118170 162302 118226
rect 162358 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 193554 118226
rect 193610 118170 193678 118226
rect 193734 118170 193802 118226
rect 193858 118170 193926 118226
rect 193982 118170 224274 118226
rect 224330 118170 224398 118226
rect 224454 118170 224522 118226
rect 224578 118170 224646 118226
rect 224702 118170 246612 118226
rect 246668 118170 246736 118226
rect 246792 118170 246860 118226
rect 246916 118170 246984 118226
rect 247040 118170 254994 118226
rect 255050 118170 255118 118226
rect 255174 118170 255242 118226
rect 255298 118170 255366 118226
rect 255422 118170 261930 118226
rect 261986 118170 262054 118226
rect 262110 118170 262178 118226
rect 262234 118170 262302 118226
rect 262358 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 346612 118226
rect 346668 118170 346736 118226
rect 346792 118170 346860 118226
rect 346916 118170 346984 118226
rect 347040 118170 361930 118226
rect 361986 118170 362054 118226
rect 362110 118170 362178 118226
rect 362234 118170 362302 118226
rect 362358 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 446612 118226
rect 446668 118170 446736 118226
rect 446792 118170 446860 118226
rect 446916 118170 446984 118226
rect 447040 118170 461930 118226
rect 461986 118170 462054 118226
rect 462110 118170 462178 118226
rect 462234 118170 462302 118226
rect 462358 118170 470034 118226
rect 470090 118170 470158 118226
rect 470214 118170 470282 118226
rect 470338 118170 470406 118226
rect 470462 118170 500754 118226
rect 500810 118170 500878 118226
rect 500934 118170 501002 118226
rect 501058 118170 501126 118226
rect 501182 118170 531474 118226
rect 531530 118170 531598 118226
rect 531654 118170 531722 118226
rect 531778 118170 531846 118226
rect 531902 118170 546612 118226
rect 546668 118170 546736 118226
rect 546792 118170 546860 118226
rect 546916 118170 546984 118226
rect 547040 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 61930 118102
rect 61986 118046 62054 118102
rect 62110 118046 62178 118102
rect 62234 118046 62302 118102
rect 62358 118046 70674 118102
rect 70730 118046 70798 118102
rect 70854 118046 70922 118102
rect 70978 118046 71046 118102
rect 71102 118046 101394 118102
rect 101450 118046 101518 118102
rect 101574 118046 101642 118102
rect 101698 118046 101766 118102
rect 101822 118046 132114 118102
rect 132170 118046 132238 118102
rect 132294 118046 132362 118102
rect 132418 118046 132486 118102
rect 132542 118046 146612 118102
rect 146668 118046 146736 118102
rect 146792 118046 146860 118102
rect 146916 118046 146984 118102
rect 147040 118046 161930 118102
rect 161986 118046 162054 118102
rect 162110 118046 162178 118102
rect 162234 118046 162302 118102
rect 162358 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 193554 118102
rect 193610 118046 193678 118102
rect 193734 118046 193802 118102
rect 193858 118046 193926 118102
rect 193982 118046 224274 118102
rect 224330 118046 224398 118102
rect 224454 118046 224522 118102
rect 224578 118046 224646 118102
rect 224702 118046 246612 118102
rect 246668 118046 246736 118102
rect 246792 118046 246860 118102
rect 246916 118046 246984 118102
rect 247040 118046 254994 118102
rect 255050 118046 255118 118102
rect 255174 118046 255242 118102
rect 255298 118046 255366 118102
rect 255422 118046 261930 118102
rect 261986 118046 262054 118102
rect 262110 118046 262178 118102
rect 262234 118046 262302 118102
rect 262358 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 346612 118102
rect 346668 118046 346736 118102
rect 346792 118046 346860 118102
rect 346916 118046 346984 118102
rect 347040 118046 361930 118102
rect 361986 118046 362054 118102
rect 362110 118046 362178 118102
rect 362234 118046 362302 118102
rect 362358 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 446612 118102
rect 446668 118046 446736 118102
rect 446792 118046 446860 118102
rect 446916 118046 446984 118102
rect 447040 118046 461930 118102
rect 461986 118046 462054 118102
rect 462110 118046 462178 118102
rect 462234 118046 462302 118102
rect 462358 118046 470034 118102
rect 470090 118046 470158 118102
rect 470214 118046 470282 118102
rect 470338 118046 470406 118102
rect 470462 118046 500754 118102
rect 500810 118046 500878 118102
rect 500934 118046 501002 118102
rect 501058 118046 501126 118102
rect 501182 118046 531474 118102
rect 531530 118046 531598 118102
rect 531654 118046 531722 118102
rect 531778 118046 531846 118102
rect 531902 118046 546612 118102
rect 546668 118046 546736 118102
rect 546792 118046 546860 118102
rect 546916 118046 546984 118102
rect 547040 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 61930 117978
rect 61986 117922 62054 117978
rect 62110 117922 62178 117978
rect 62234 117922 62302 117978
rect 62358 117922 70674 117978
rect 70730 117922 70798 117978
rect 70854 117922 70922 117978
rect 70978 117922 71046 117978
rect 71102 117922 101394 117978
rect 101450 117922 101518 117978
rect 101574 117922 101642 117978
rect 101698 117922 101766 117978
rect 101822 117922 132114 117978
rect 132170 117922 132238 117978
rect 132294 117922 132362 117978
rect 132418 117922 132486 117978
rect 132542 117922 146612 117978
rect 146668 117922 146736 117978
rect 146792 117922 146860 117978
rect 146916 117922 146984 117978
rect 147040 117922 161930 117978
rect 161986 117922 162054 117978
rect 162110 117922 162178 117978
rect 162234 117922 162302 117978
rect 162358 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 193554 117978
rect 193610 117922 193678 117978
rect 193734 117922 193802 117978
rect 193858 117922 193926 117978
rect 193982 117922 224274 117978
rect 224330 117922 224398 117978
rect 224454 117922 224522 117978
rect 224578 117922 224646 117978
rect 224702 117922 246612 117978
rect 246668 117922 246736 117978
rect 246792 117922 246860 117978
rect 246916 117922 246984 117978
rect 247040 117922 254994 117978
rect 255050 117922 255118 117978
rect 255174 117922 255242 117978
rect 255298 117922 255366 117978
rect 255422 117922 261930 117978
rect 261986 117922 262054 117978
rect 262110 117922 262178 117978
rect 262234 117922 262302 117978
rect 262358 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 346612 117978
rect 346668 117922 346736 117978
rect 346792 117922 346860 117978
rect 346916 117922 346984 117978
rect 347040 117922 361930 117978
rect 361986 117922 362054 117978
rect 362110 117922 362178 117978
rect 362234 117922 362302 117978
rect 362358 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 446612 117978
rect 446668 117922 446736 117978
rect 446792 117922 446860 117978
rect 446916 117922 446984 117978
rect 447040 117922 461930 117978
rect 461986 117922 462054 117978
rect 462110 117922 462178 117978
rect 462234 117922 462302 117978
rect 462358 117922 470034 117978
rect 470090 117922 470158 117978
rect 470214 117922 470282 117978
rect 470338 117922 470406 117978
rect 470462 117922 500754 117978
rect 500810 117922 500878 117978
rect 500934 117922 501002 117978
rect 501058 117922 501126 117978
rect 501182 117922 531474 117978
rect 531530 117922 531598 117978
rect 531654 117922 531722 117978
rect 531778 117922 531846 117978
rect 531902 117922 546612 117978
rect 546668 117922 546736 117978
rect 546792 117922 546860 117978
rect 546916 117922 546984 117978
rect 547040 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 61130 112350
rect 61186 112294 61254 112350
rect 61310 112294 61378 112350
rect 61434 112294 61502 112350
rect 61558 112294 66954 112350
rect 67010 112294 67078 112350
rect 67134 112294 67202 112350
rect 67258 112294 67326 112350
rect 67382 112294 97674 112350
rect 97730 112294 97798 112350
rect 97854 112294 97922 112350
rect 97978 112294 98046 112350
rect 98102 112294 128394 112350
rect 128450 112294 128518 112350
rect 128574 112294 128642 112350
rect 128698 112294 128766 112350
rect 128822 112294 145812 112350
rect 145868 112294 145936 112350
rect 145992 112294 146060 112350
rect 146116 112294 146184 112350
rect 146240 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 161130 112350
rect 161186 112294 161254 112350
rect 161310 112294 161378 112350
rect 161434 112294 161502 112350
rect 161558 112294 189834 112350
rect 189890 112294 189958 112350
rect 190014 112294 190082 112350
rect 190138 112294 190206 112350
rect 190262 112294 220554 112350
rect 220610 112294 220678 112350
rect 220734 112294 220802 112350
rect 220858 112294 220926 112350
rect 220982 112294 245812 112350
rect 245868 112294 245936 112350
rect 245992 112294 246060 112350
rect 246116 112294 246184 112350
rect 246240 112294 251274 112350
rect 251330 112294 251398 112350
rect 251454 112294 251522 112350
rect 251578 112294 251646 112350
rect 251702 112294 261130 112350
rect 261186 112294 261254 112350
rect 261310 112294 261378 112350
rect 261434 112294 261502 112350
rect 261558 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 345812 112350
rect 345868 112294 345936 112350
rect 345992 112294 346060 112350
rect 346116 112294 346184 112350
rect 346240 112294 361130 112350
rect 361186 112294 361254 112350
rect 361310 112294 361378 112350
rect 361434 112294 361502 112350
rect 361558 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 445812 112350
rect 445868 112294 445936 112350
rect 445992 112294 446060 112350
rect 446116 112294 446184 112350
rect 446240 112294 461130 112350
rect 461186 112294 461254 112350
rect 461310 112294 461378 112350
rect 461434 112294 461502 112350
rect 461558 112294 466314 112350
rect 466370 112294 466438 112350
rect 466494 112294 466562 112350
rect 466618 112294 466686 112350
rect 466742 112294 497034 112350
rect 497090 112294 497158 112350
rect 497214 112294 497282 112350
rect 497338 112294 497406 112350
rect 497462 112294 527754 112350
rect 527810 112294 527878 112350
rect 527934 112294 528002 112350
rect 528058 112294 528126 112350
rect 528182 112294 545812 112350
rect 545868 112294 545936 112350
rect 545992 112294 546060 112350
rect 546116 112294 546184 112350
rect 546240 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 61130 112226
rect 61186 112170 61254 112226
rect 61310 112170 61378 112226
rect 61434 112170 61502 112226
rect 61558 112170 66954 112226
rect 67010 112170 67078 112226
rect 67134 112170 67202 112226
rect 67258 112170 67326 112226
rect 67382 112170 97674 112226
rect 97730 112170 97798 112226
rect 97854 112170 97922 112226
rect 97978 112170 98046 112226
rect 98102 112170 128394 112226
rect 128450 112170 128518 112226
rect 128574 112170 128642 112226
rect 128698 112170 128766 112226
rect 128822 112170 145812 112226
rect 145868 112170 145936 112226
rect 145992 112170 146060 112226
rect 146116 112170 146184 112226
rect 146240 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 161130 112226
rect 161186 112170 161254 112226
rect 161310 112170 161378 112226
rect 161434 112170 161502 112226
rect 161558 112170 189834 112226
rect 189890 112170 189958 112226
rect 190014 112170 190082 112226
rect 190138 112170 190206 112226
rect 190262 112170 220554 112226
rect 220610 112170 220678 112226
rect 220734 112170 220802 112226
rect 220858 112170 220926 112226
rect 220982 112170 245812 112226
rect 245868 112170 245936 112226
rect 245992 112170 246060 112226
rect 246116 112170 246184 112226
rect 246240 112170 251274 112226
rect 251330 112170 251398 112226
rect 251454 112170 251522 112226
rect 251578 112170 251646 112226
rect 251702 112170 261130 112226
rect 261186 112170 261254 112226
rect 261310 112170 261378 112226
rect 261434 112170 261502 112226
rect 261558 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 345812 112226
rect 345868 112170 345936 112226
rect 345992 112170 346060 112226
rect 346116 112170 346184 112226
rect 346240 112170 361130 112226
rect 361186 112170 361254 112226
rect 361310 112170 361378 112226
rect 361434 112170 361502 112226
rect 361558 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 445812 112226
rect 445868 112170 445936 112226
rect 445992 112170 446060 112226
rect 446116 112170 446184 112226
rect 446240 112170 461130 112226
rect 461186 112170 461254 112226
rect 461310 112170 461378 112226
rect 461434 112170 461502 112226
rect 461558 112170 466314 112226
rect 466370 112170 466438 112226
rect 466494 112170 466562 112226
rect 466618 112170 466686 112226
rect 466742 112170 497034 112226
rect 497090 112170 497158 112226
rect 497214 112170 497282 112226
rect 497338 112170 497406 112226
rect 497462 112170 527754 112226
rect 527810 112170 527878 112226
rect 527934 112170 528002 112226
rect 528058 112170 528126 112226
rect 528182 112170 545812 112226
rect 545868 112170 545936 112226
rect 545992 112170 546060 112226
rect 546116 112170 546184 112226
rect 546240 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 61130 112102
rect 61186 112046 61254 112102
rect 61310 112046 61378 112102
rect 61434 112046 61502 112102
rect 61558 112046 66954 112102
rect 67010 112046 67078 112102
rect 67134 112046 67202 112102
rect 67258 112046 67326 112102
rect 67382 112046 97674 112102
rect 97730 112046 97798 112102
rect 97854 112046 97922 112102
rect 97978 112046 98046 112102
rect 98102 112046 128394 112102
rect 128450 112046 128518 112102
rect 128574 112046 128642 112102
rect 128698 112046 128766 112102
rect 128822 112046 145812 112102
rect 145868 112046 145936 112102
rect 145992 112046 146060 112102
rect 146116 112046 146184 112102
rect 146240 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 161130 112102
rect 161186 112046 161254 112102
rect 161310 112046 161378 112102
rect 161434 112046 161502 112102
rect 161558 112046 189834 112102
rect 189890 112046 189958 112102
rect 190014 112046 190082 112102
rect 190138 112046 190206 112102
rect 190262 112046 220554 112102
rect 220610 112046 220678 112102
rect 220734 112046 220802 112102
rect 220858 112046 220926 112102
rect 220982 112046 245812 112102
rect 245868 112046 245936 112102
rect 245992 112046 246060 112102
rect 246116 112046 246184 112102
rect 246240 112046 251274 112102
rect 251330 112046 251398 112102
rect 251454 112046 251522 112102
rect 251578 112046 251646 112102
rect 251702 112046 261130 112102
rect 261186 112046 261254 112102
rect 261310 112046 261378 112102
rect 261434 112046 261502 112102
rect 261558 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 345812 112102
rect 345868 112046 345936 112102
rect 345992 112046 346060 112102
rect 346116 112046 346184 112102
rect 346240 112046 361130 112102
rect 361186 112046 361254 112102
rect 361310 112046 361378 112102
rect 361434 112046 361502 112102
rect 361558 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 445812 112102
rect 445868 112046 445936 112102
rect 445992 112046 446060 112102
rect 446116 112046 446184 112102
rect 446240 112046 461130 112102
rect 461186 112046 461254 112102
rect 461310 112046 461378 112102
rect 461434 112046 461502 112102
rect 461558 112046 466314 112102
rect 466370 112046 466438 112102
rect 466494 112046 466562 112102
rect 466618 112046 466686 112102
rect 466742 112046 497034 112102
rect 497090 112046 497158 112102
rect 497214 112046 497282 112102
rect 497338 112046 497406 112102
rect 497462 112046 527754 112102
rect 527810 112046 527878 112102
rect 527934 112046 528002 112102
rect 528058 112046 528126 112102
rect 528182 112046 545812 112102
rect 545868 112046 545936 112102
rect 545992 112046 546060 112102
rect 546116 112046 546184 112102
rect 546240 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 61130 111978
rect 61186 111922 61254 111978
rect 61310 111922 61378 111978
rect 61434 111922 61502 111978
rect 61558 111922 66954 111978
rect 67010 111922 67078 111978
rect 67134 111922 67202 111978
rect 67258 111922 67326 111978
rect 67382 111922 97674 111978
rect 97730 111922 97798 111978
rect 97854 111922 97922 111978
rect 97978 111922 98046 111978
rect 98102 111922 128394 111978
rect 128450 111922 128518 111978
rect 128574 111922 128642 111978
rect 128698 111922 128766 111978
rect 128822 111922 145812 111978
rect 145868 111922 145936 111978
rect 145992 111922 146060 111978
rect 146116 111922 146184 111978
rect 146240 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 161130 111978
rect 161186 111922 161254 111978
rect 161310 111922 161378 111978
rect 161434 111922 161502 111978
rect 161558 111922 189834 111978
rect 189890 111922 189958 111978
rect 190014 111922 190082 111978
rect 190138 111922 190206 111978
rect 190262 111922 220554 111978
rect 220610 111922 220678 111978
rect 220734 111922 220802 111978
rect 220858 111922 220926 111978
rect 220982 111922 245812 111978
rect 245868 111922 245936 111978
rect 245992 111922 246060 111978
rect 246116 111922 246184 111978
rect 246240 111922 251274 111978
rect 251330 111922 251398 111978
rect 251454 111922 251522 111978
rect 251578 111922 251646 111978
rect 251702 111922 261130 111978
rect 261186 111922 261254 111978
rect 261310 111922 261378 111978
rect 261434 111922 261502 111978
rect 261558 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 345812 111978
rect 345868 111922 345936 111978
rect 345992 111922 346060 111978
rect 346116 111922 346184 111978
rect 346240 111922 361130 111978
rect 361186 111922 361254 111978
rect 361310 111922 361378 111978
rect 361434 111922 361502 111978
rect 361558 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 445812 111978
rect 445868 111922 445936 111978
rect 445992 111922 446060 111978
rect 446116 111922 446184 111978
rect 446240 111922 461130 111978
rect 461186 111922 461254 111978
rect 461310 111922 461378 111978
rect 461434 111922 461502 111978
rect 461558 111922 466314 111978
rect 466370 111922 466438 111978
rect 466494 111922 466562 111978
rect 466618 111922 466686 111978
rect 466742 111922 497034 111978
rect 497090 111922 497158 111978
rect 497214 111922 497282 111978
rect 497338 111922 497406 111978
rect 497462 111922 527754 111978
rect 527810 111922 527878 111978
rect 527934 111922 528002 111978
rect 528058 111922 528126 111978
rect 528182 111922 545812 111978
rect 545868 111922 545936 111978
rect 545992 111922 546060 111978
rect 546116 111922 546184 111978
rect 546240 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 61930 100350
rect 61986 100294 62054 100350
rect 62110 100294 62178 100350
rect 62234 100294 62302 100350
rect 62358 100294 70674 100350
rect 70730 100294 70798 100350
rect 70854 100294 70922 100350
rect 70978 100294 71046 100350
rect 71102 100294 101394 100350
rect 101450 100294 101518 100350
rect 101574 100294 101642 100350
rect 101698 100294 101766 100350
rect 101822 100294 132114 100350
rect 132170 100294 132238 100350
rect 132294 100294 132362 100350
rect 132418 100294 132486 100350
rect 132542 100294 146612 100350
rect 146668 100294 146736 100350
rect 146792 100294 146860 100350
rect 146916 100294 146984 100350
rect 147040 100294 161930 100350
rect 161986 100294 162054 100350
rect 162110 100294 162178 100350
rect 162234 100294 162302 100350
rect 162358 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 193554 100350
rect 193610 100294 193678 100350
rect 193734 100294 193802 100350
rect 193858 100294 193926 100350
rect 193982 100294 224274 100350
rect 224330 100294 224398 100350
rect 224454 100294 224522 100350
rect 224578 100294 224646 100350
rect 224702 100294 246612 100350
rect 246668 100294 246736 100350
rect 246792 100294 246860 100350
rect 246916 100294 246984 100350
rect 247040 100294 254994 100350
rect 255050 100294 255118 100350
rect 255174 100294 255242 100350
rect 255298 100294 255366 100350
rect 255422 100294 261930 100350
rect 261986 100294 262054 100350
rect 262110 100294 262178 100350
rect 262234 100294 262302 100350
rect 262358 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 346612 100350
rect 346668 100294 346736 100350
rect 346792 100294 346860 100350
rect 346916 100294 346984 100350
rect 347040 100294 361930 100350
rect 361986 100294 362054 100350
rect 362110 100294 362178 100350
rect 362234 100294 362302 100350
rect 362358 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 446612 100350
rect 446668 100294 446736 100350
rect 446792 100294 446860 100350
rect 446916 100294 446984 100350
rect 447040 100294 461930 100350
rect 461986 100294 462054 100350
rect 462110 100294 462178 100350
rect 462234 100294 462302 100350
rect 462358 100294 470034 100350
rect 470090 100294 470158 100350
rect 470214 100294 470282 100350
rect 470338 100294 470406 100350
rect 470462 100294 500754 100350
rect 500810 100294 500878 100350
rect 500934 100294 501002 100350
rect 501058 100294 501126 100350
rect 501182 100294 531474 100350
rect 531530 100294 531598 100350
rect 531654 100294 531722 100350
rect 531778 100294 531846 100350
rect 531902 100294 546612 100350
rect 546668 100294 546736 100350
rect 546792 100294 546860 100350
rect 546916 100294 546984 100350
rect 547040 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 61930 100226
rect 61986 100170 62054 100226
rect 62110 100170 62178 100226
rect 62234 100170 62302 100226
rect 62358 100170 70674 100226
rect 70730 100170 70798 100226
rect 70854 100170 70922 100226
rect 70978 100170 71046 100226
rect 71102 100170 101394 100226
rect 101450 100170 101518 100226
rect 101574 100170 101642 100226
rect 101698 100170 101766 100226
rect 101822 100170 132114 100226
rect 132170 100170 132238 100226
rect 132294 100170 132362 100226
rect 132418 100170 132486 100226
rect 132542 100170 146612 100226
rect 146668 100170 146736 100226
rect 146792 100170 146860 100226
rect 146916 100170 146984 100226
rect 147040 100170 161930 100226
rect 161986 100170 162054 100226
rect 162110 100170 162178 100226
rect 162234 100170 162302 100226
rect 162358 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 193554 100226
rect 193610 100170 193678 100226
rect 193734 100170 193802 100226
rect 193858 100170 193926 100226
rect 193982 100170 224274 100226
rect 224330 100170 224398 100226
rect 224454 100170 224522 100226
rect 224578 100170 224646 100226
rect 224702 100170 246612 100226
rect 246668 100170 246736 100226
rect 246792 100170 246860 100226
rect 246916 100170 246984 100226
rect 247040 100170 254994 100226
rect 255050 100170 255118 100226
rect 255174 100170 255242 100226
rect 255298 100170 255366 100226
rect 255422 100170 261930 100226
rect 261986 100170 262054 100226
rect 262110 100170 262178 100226
rect 262234 100170 262302 100226
rect 262358 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 346612 100226
rect 346668 100170 346736 100226
rect 346792 100170 346860 100226
rect 346916 100170 346984 100226
rect 347040 100170 361930 100226
rect 361986 100170 362054 100226
rect 362110 100170 362178 100226
rect 362234 100170 362302 100226
rect 362358 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 446612 100226
rect 446668 100170 446736 100226
rect 446792 100170 446860 100226
rect 446916 100170 446984 100226
rect 447040 100170 461930 100226
rect 461986 100170 462054 100226
rect 462110 100170 462178 100226
rect 462234 100170 462302 100226
rect 462358 100170 470034 100226
rect 470090 100170 470158 100226
rect 470214 100170 470282 100226
rect 470338 100170 470406 100226
rect 470462 100170 500754 100226
rect 500810 100170 500878 100226
rect 500934 100170 501002 100226
rect 501058 100170 501126 100226
rect 501182 100170 531474 100226
rect 531530 100170 531598 100226
rect 531654 100170 531722 100226
rect 531778 100170 531846 100226
rect 531902 100170 546612 100226
rect 546668 100170 546736 100226
rect 546792 100170 546860 100226
rect 546916 100170 546984 100226
rect 547040 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 61930 100102
rect 61986 100046 62054 100102
rect 62110 100046 62178 100102
rect 62234 100046 62302 100102
rect 62358 100046 70674 100102
rect 70730 100046 70798 100102
rect 70854 100046 70922 100102
rect 70978 100046 71046 100102
rect 71102 100046 101394 100102
rect 101450 100046 101518 100102
rect 101574 100046 101642 100102
rect 101698 100046 101766 100102
rect 101822 100046 132114 100102
rect 132170 100046 132238 100102
rect 132294 100046 132362 100102
rect 132418 100046 132486 100102
rect 132542 100046 146612 100102
rect 146668 100046 146736 100102
rect 146792 100046 146860 100102
rect 146916 100046 146984 100102
rect 147040 100046 161930 100102
rect 161986 100046 162054 100102
rect 162110 100046 162178 100102
rect 162234 100046 162302 100102
rect 162358 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 193554 100102
rect 193610 100046 193678 100102
rect 193734 100046 193802 100102
rect 193858 100046 193926 100102
rect 193982 100046 224274 100102
rect 224330 100046 224398 100102
rect 224454 100046 224522 100102
rect 224578 100046 224646 100102
rect 224702 100046 246612 100102
rect 246668 100046 246736 100102
rect 246792 100046 246860 100102
rect 246916 100046 246984 100102
rect 247040 100046 254994 100102
rect 255050 100046 255118 100102
rect 255174 100046 255242 100102
rect 255298 100046 255366 100102
rect 255422 100046 261930 100102
rect 261986 100046 262054 100102
rect 262110 100046 262178 100102
rect 262234 100046 262302 100102
rect 262358 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 346612 100102
rect 346668 100046 346736 100102
rect 346792 100046 346860 100102
rect 346916 100046 346984 100102
rect 347040 100046 361930 100102
rect 361986 100046 362054 100102
rect 362110 100046 362178 100102
rect 362234 100046 362302 100102
rect 362358 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 446612 100102
rect 446668 100046 446736 100102
rect 446792 100046 446860 100102
rect 446916 100046 446984 100102
rect 447040 100046 461930 100102
rect 461986 100046 462054 100102
rect 462110 100046 462178 100102
rect 462234 100046 462302 100102
rect 462358 100046 470034 100102
rect 470090 100046 470158 100102
rect 470214 100046 470282 100102
rect 470338 100046 470406 100102
rect 470462 100046 500754 100102
rect 500810 100046 500878 100102
rect 500934 100046 501002 100102
rect 501058 100046 501126 100102
rect 501182 100046 531474 100102
rect 531530 100046 531598 100102
rect 531654 100046 531722 100102
rect 531778 100046 531846 100102
rect 531902 100046 546612 100102
rect 546668 100046 546736 100102
rect 546792 100046 546860 100102
rect 546916 100046 546984 100102
rect 547040 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 61930 99978
rect 61986 99922 62054 99978
rect 62110 99922 62178 99978
rect 62234 99922 62302 99978
rect 62358 99922 70674 99978
rect 70730 99922 70798 99978
rect 70854 99922 70922 99978
rect 70978 99922 71046 99978
rect 71102 99922 101394 99978
rect 101450 99922 101518 99978
rect 101574 99922 101642 99978
rect 101698 99922 101766 99978
rect 101822 99922 132114 99978
rect 132170 99922 132238 99978
rect 132294 99922 132362 99978
rect 132418 99922 132486 99978
rect 132542 99922 146612 99978
rect 146668 99922 146736 99978
rect 146792 99922 146860 99978
rect 146916 99922 146984 99978
rect 147040 99922 161930 99978
rect 161986 99922 162054 99978
rect 162110 99922 162178 99978
rect 162234 99922 162302 99978
rect 162358 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 193554 99978
rect 193610 99922 193678 99978
rect 193734 99922 193802 99978
rect 193858 99922 193926 99978
rect 193982 99922 224274 99978
rect 224330 99922 224398 99978
rect 224454 99922 224522 99978
rect 224578 99922 224646 99978
rect 224702 99922 246612 99978
rect 246668 99922 246736 99978
rect 246792 99922 246860 99978
rect 246916 99922 246984 99978
rect 247040 99922 254994 99978
rect 255050 99922 255118 99978
rect 255174 99922 255242 99978
rect 255298 99922 255366 99978
rect 255422 99922 261930 99978
rect 261986 99922 262054 99978
rect 262110 99922 262178 99978
rect 262234 99922 262302 99978
rect 262358 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 346612 99978
rect 346668 99922 346736 99978
rect 346792 99922 346860 99978
rect 346916 99922 346984 99978
rect 347040 99922 361930 99978
rect 361986 99922 362054 99978
rect 362110 99922 362178 99978
rect 362234 99922 362302 99978
rect 362358 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 446612 99978
rect 446668 99922 446736 99978
rect 446792 99922 446860 99978
rect 446916 99922 446984 99978
rect 447040 99922 461930 99978
rect 461986 99922 462054 99978
rect 462110 99922 462178 99978
rect 462234 99922 462302 99978
rect 462358 99922 470034 99978
rect 470090 99922 470158 99978
rect 470214 99922 470282 99978
rect 470338 99922 470406 99978
rect 470462 99922 500754 99978
rect 500810 99922 500878 99978
rect 500934 99922 501002 99978
rect 501058 99922 501126 99978
rect 501182 99922 531474 99978
rect 531530 99922 531598 99978
rect 531654 99922 531722 99978
rect 531778 99922 531846 99978
rect 531902 99922 546612 99978
rect 546668 99922 546736 99978
rect 546792 99922 546860 99978
rect 546916 99922 546984 99978
rect 547040 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 61130 94350
rect 61186 94294 61254 94350
rect 61310 94294 61378 94350
rect 61434 94294 61502 94350
rect 61558 94294 66954 94350
rect 67010 94294 67078 94350
rect 67134 94294 67202 94350
rect 67258 94294 67326 94350
rect 67382 94294 97674 94350
rect 97730 94294 97798 94350
rect 97854 94294 97922 94350
rect 97978 94294 98046 94350
rect 98102 94294 128394 94350
rect 128450 94294 128518 94350
rect 128574 94294 128642 94350
rect 128698 94294 128766 94350
rect 128822 94294 145812 94350
rect 145868 94294 145936 94350
rect 145992 94294 146060 94350
rect 146116 94294 146184 94350
rect 146240 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 161130 94350
rect 161186 94294 161254 94350
rect 161310 94294 161378 94350
rect 161434 94294 161502 94350
rect 161558 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 245812 94350
rect 245868 94294 245936 94350
rect 245992 94294 246060 94350
rect 246116 94294 246184 94350
rect 246240 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 261130 94350
rect 261186 94294 261254 94350
rect 261310 94294 261378 94350
rect 261434 94294 261502 94350
rect 261558 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 345812 94350
rect 345868 94294 345936 94350
rect 345992 94294 346060 94350
rect 346116 94294 346184 94350
rect 346240 94294 361130 94350
rect 361186 94294 361254 94350
rect 361310 94294 361378 94350
rect 361434 94294 361502 94350
rect 361558 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 404874 94350
rect 404930 94294 404998 94350
rect 405054 94294 405122 94350
rect 405178 94294 405246 94350
rect 405302 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 445812 94350
rect 445868 94294 445936 94350
rect 445992 94294 446060 94350
rect 446116 94294 446184 94350
rect 446240 94294 461130 94350
rect 461186 94294 461254 94350
rect 461310 94294 461378 94350
rect 461434 94294 461502 94350
rect 461558 94294 466314 94350
rect 466370 94294 466438 94350
rect 466494 94294 466562 94350
rect 466618 94294 466686 94350
rect 466742 94294 497034 94350
rect 497090 94294 497158 94350
rect 497214 94294 497282 94350
rect 497338 94294 497406 94350
rect 497462 94294 527754 94350
rect 527810 94294 527878 94350
rect 527934 94294 528002 94350
rect 528058 94294 528126 94350
rect 528182 94294 545812 94350
rect 545868 94294 545936 94350
rect 545992 94294 546060 94350
rect 546116 94294 546184 94350
rect 546240 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 61130 94226
rect 61186 94170 61254 94226
rect 61310 94170 61378 94226
rect 61434 94170 61502 94226
rect 61558 94170 66954 94226
rect 67010 94170 67078 94226
rect 67134 94170 67202 94226
rect 67258 94170 67326 94226
rect 67382 94170 97674 94226
rect 97730 94170 97798 94226
rect 97854 94170 97922 94226
rect 97978 94170 98046 94226
rect 98102 94170 128394 94226
rect 128450 94170 128518 94226
rect 128574 94170 128642 94226
rect 128698 94170 128766 94226
rect 128822 94170 145812 94226
rect 145868 94170 145936 94226
rect 145992 94170 146060 94226
rect 146116 94170 146184 94226
rect 146240 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 161130 94226
rect 161186 94170 161254 94226
rect 161310 94170 161378 94226
rect 161434 94170 161502 94226
rect 161558 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 245812 94226
rect 245868 94170 245936 94226
rect 245992 94170 246060 94226
rect 246116 94170 246184 94226
rect 246240 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 261130 94226
rect 261186 94170 261254 94226
rect 261310 94170 261378 94226
rect 261434 94170 261502 94226
rect 261558 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 345812 94226
rect 345868 94170 345936 94226
rect 345992 94170 346060 94226
rect 346116 94170 346184 94226
rect 346240 94170 361130 94226
rect 361186 94170 361254 94226
rect 361310 94170 361378 94226
rect 361434 94170 361502 94226
rect 361558 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 404874 94226
rect 404930 94170 404998 94226
rect 405054 94170 405122 94226
rect 405178 94170 405246 94226
rect 405302 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 445812 94226
rect 445868 94170 445936 94226
rect 445992 94170 446060 94226
rect 446116 94170 446184 94226
rect 446240 94170 461130 94226
rect 461186 94170 461254 94226
rect 461310 94170 461378 94226
rect 461434 94170 461502 94226
rect 461558 94170 466314 94226
rect 466370 94170 466438 94226
rect 466494 94170 466562 94226
rect 466618 94170 466686 94226
rect 466742 94170 497034 94226
rect 497090 94170 497158 94226
rect 497214 94170 497282 94226
rect 497338 94170 497406 94226
rect 497462 94170 527754 94226
rect 527810 94170 527878 94226
rect 527934 94170 528002 94226
rect 528058 94170 528126 94226
rect 528182 94170 545812 94226
rect 545868 94170 545936 94226
rect 545992 94170 546060 94226
rect 546116 94170 546184 94226
rect 546240 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 61130 94102
rect 61186 94046 61254 94102
rect 61310 94046 61378 94102
rect 61434 94046 61502 94102
rect 61558 94046 66954 94102
rect 67010 94046 67078 94102
rect 67134 94046 67202 94102
rect 67258 94046 67326 94102
rect 67382 94046 97674 94102
rect 97730 94046 97798 94102
rect 97854 94046 97922 94102
rect 97978 94046 98046 94102
rect 98102 94046 128394 94102
rect 128450 94046 128518 94102
rect 128574 94046 128642 94102
rect 128698 94046 128766 94102
rect 128822 94046 145812 94102
rect 145868 94046 145936 94102
rect 145992 94046 146060 94102
rect 146116 94046 146184 94102
rect 146240 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 161130 94102
rect 161186 94046 161254 94102
rect 161310 94046 161378 94102
rect 161434 94046 161502 94102
rect 161558 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 245812 94102
rect 245868 94046 245936 94102
rect 245992 94046 246060 94102
rect 246116 94046 246184 94102
rect 246240 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 261130 94102
rect 261186 94046 261254 94102
rect 261310 94046 261378 94102
rect 261434 94046 261502 94102
rect 261558 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 345812 94102
rect 345868 94046 345936 94102
rect 345992 94046 346060 94102
rect 346116 94046 346184 94102
rect 346240 94046 361130 94102
rect 361186 94046 361254 94102
rect 361310 94046 361378 94102
rect 361434 94046 361502 94102
rect 361558 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 404874 94102
rect 404930 94046 404998 94102
rect 405054 94046 405122 94102
rect 405178 94046 405246 94102
rect 405302 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 445812 94102
rect 445868 94046 445936 94102
rect 445992 94046 446060 94102
rect 446116 94046 446184 94102
rect 446240 94046 461130 94102
rect 461186 94046 461254 94102
rect 461310 94046 461378 94102
rect 461434 94046 461502 94102
rect 461558 94046 466314 94102
rect 466370 94046 466438 94102
rect 466494 94046 466562 94102
rect 466618 94046 466686 94102
rect 466742 94046 497034 94102
rect 497090 94046 497158 94102
rect 497214 94046 497282 94102
rect 497338 94046 497406 94102
rect 497462 94046 527754 94102
rect 527810 94046 527878 94102
rect 527934 94046 528002 94102
rect 528058 94046 528126 94102
rect 528182 94046 545812 94102
rect 545868 94046 545936 94102
rect 545992 94046 546060 94102
rect 546116 94046 546184 94102
rect 546240 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 61130 93978
rect 61186 93922 61254 93978
rect 61310 93922 61378 93978
rect 61434 93922 61502 93978
rect 61558 93922 66954 93978
rect 67010 93922 67078 93978
rect 67134 93922 67202 93978
rect 67258 93922 67326 93978
rect 67382 93922 97674 93978
rect 97730 93922 97798 93978
rect 97854 93922 97922 93978
rect 97978 93922 98046 93978
rect 98102 93922 128394 93978
rect 128450 93922 128518 93978
rect 128574 93922 128642 93978
rect 128698 93922 128766 93978
rect 128822 93922 145812 93978
rect 145868 93922 145936 93978
rect 145992 93922 146060 93978
rect 146116 93922 146184 93978
rect 146240 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 161130 93978
rect 161186 93922 161254 93978
rect 161310 93922 161378 93978
rect 161434 93922 161502 93978
rect 161558 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 245812 93978
rect 245868 93922 245936 93978
rect 245992 93922 246060 93978
rect 246116 93922 246184 93978
rect 246240 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 261130 93978
rect 261186 93922 261254 93978
rect 261310 93922 261378 93978
rect 261434 93922 261502 93978
rect 261558 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 345812 93978
rect 345868 93922 345936 93978
rect 345992 93922 346060 93978
rect 346116 93922 346184 93978
rect 346240 93922 361130 93978
rect 361186 93922 361254 93978
rect 361310 93922 361378 93978
rect 361434 93922 361502 93978
rect 361558 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 404874 93978
rect 404930 93922 404998 93978
rect 405054 93922 405122 93978
rect 405178 93922 405246 93978
rect 405302 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 445812 93978
rect 445868 93922 445936 93978
rect 445992 93922 446060 93978
rect 446116 93922 446184 93978
rect 446240 93922 461130 93978
rect 461186 93922 461254 93978
rect 461310 93922 461378 93978
rect 461434 93922 461502 93978
rect 461558 93922 466314 93978
rect 466370 93922 466438 93978
rect 466494 93922 466562 93978
rect 466618 93922 466686 93978
rect 466742 93922 497034 93978
rect 497090 93922 497158 93978
rect 497214 93922 497282 93978
rect 497338 93922 497406 93978
rect 497462 93922 527754 93978
rect 527810 93922 527878 93978
rect 527934 93922 528002 93978
rect 528058 93922 528126 93978
rect 528182 93922 545812 93978
rect 545868 93922 545936 93978
rect 545992 93922 546060 93978
rect 546116 93922 546184 93978
rect 546240 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 61930 82350
rect 61986 82294 62054 82350
rect 62110 82294 62178 82350
rect 62234 82294 62302 82350
rect 62358 82294 70674 82350
rect 70730 82294 70798 82350
rect 70854 82294 70922 82350
rect 70978 82294 71046 82350
rect 71102 82294 101394 82350
rect 101450 82294 101518 82350
rect 101574 82294 101642 82350
rect 101698 82294 101766 82350
rect 101822 82294 132114 82350
rect 132170 82294 132238 82350
rect 132294 82294 132362 82350
rect 132418 82294 132486 82350
rect 132542 82294 146612 82350
rect 146668 82294 146736 82350
rect 146792 82294 146860 82350
rect 146916 82294 146984 82350
rect 147040 82294 161930 82350
rect 161986 82294 162054 82350
rect 162110 82294 162178 82350
rect 162234 82294 162302 82350
rect 162358 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 224274 82350
rect 224330 82294 224398 82350
rect 224454 82294 224522 82350
rect 224578 82294 224646 82350
rect 224702 82294 246612 82350
rect 246668 82294 246736 82350
rect 246792 82294 246860 82350
rect 246916 82294 246984 82350
rect 247040 82294 254994 82350
rect 255050 82294 255118 82350
rect 255174 82294 255242 82350
rect 255298 82294 255366 82350
rect 255422 82294 261930 82350
rect 261986 82294 262054 82350
rect 262110 82294 262178 82350
rect 262234 82294 262302 82350
rect 262358 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 316434 82350
rect 316490 82294 316558 82350
rect 316614 82294 316682 82350
rect 316738 82294 316806 82350
rect 316862 82294 346612 82350
rect 346668 82294 346736 82350
rect 346792 82294 346860 82350
rect 346916 82294 346984 82350
rect 347040 82294 361930 82350
rect 361986 82294 362054 82350
rect 362110 82294 362178 82350
rect 362234 82294 362302 82350
rect 362358 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 408594 82350
rect 408650 82294 408718 82350
rect 408774 82294 408842 82350
rect 408898 82294 408966 82350
rect 409022 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 446612 82350
rect 446668 82294 446736 82350
rect 446792 82294 446860 82350
rect 446916 82294 446984 82350
rect 447040 82294 461930 82350
rect 461986 82294 462054 82350
rect 462110 82294 462178 82350
rect 462234 82294 462302 82350
rect 462358 82294 470034 82350
rect 470090 82294 470158 82350
rect 470214 82294 470282 82350
rect 470338 82294 470406 82350
rect 470462 82294 500754 82350
rect 500810 82294 500878 82350
rect 500934 82294 501002 82350
rect 501058 82294 501126 82350
rect 501182 82294 531474 82350
rect 531530 82294 531598 82350
rect 531654 82294 531722 82350
rect 531778 82294 531846 82350
rect 531902 82294 546612 82350
rect 546668 82294 546736 82350
rect 546792 82294 546860 82350
rect 546916 82294 546984 82350
rect 547040 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 61930 82226
rect 61986 82170 62054 82226
rect 62110 82170 62178 82226
rect 62234 82170 62302 82226
rect 62358 82170 70674 82226
rect 70730 82170 70798 82226
rect 70854 82170 70922 82226
rect 70978 82170 71046 82226
rect 71102 82170 101394 82226
rect 101450 82170 101518 82226
rect 101574 82170 101642 82226
rect 101698 82170 101766 82226
rect 101822 82170 132114 82226
rect 132170 82170 132238 82226
rect 132294 82170 132362 82226
rect 132418 82170 132486 82226
rect 132542 82170 146612 82226
rect 146668 82170 146736 82226
rect 146792 82170 146860 82226
rect 146916 82170 146984 82226
rect 147040 82170 161930 82226
rect 161986 82170 162054 82226
rect 162110 82170 162178 82226
rect 162234 82170 162302 82226
rect 162358 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 224274 82226
rect 224330 82170 224398 82226
rect 224454 82170 224522 82226
rect 224578 82170 224646 82226
rect 224702 82170 246612 82226
rect 246668 82170 246736 82226
rect 246792 82170 246860 82226
rect 246916 82170 246984 82226
rect 247040 82170 254994 82226
rect 255050 82170 255118 82226
rect 255174 82170 255242 82226
rect 255298 82170 255366 82226
rect 255422 82170 261930 82226
rect 261986 82170 262054 82226
rect 262110 82170 262178 82226
rect 262234 82170 262302 82226
rect 262358 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 316434 82226
rect 316490 82170 316558 82226
rect 316614 82170 316682 82226
rect 316738 82170 316806 82226
rect 316862 82170 346612 82226
rect 346668 82170 346736 82226
rect 346792 82170 346860 82226
rect 346916 82170 346984 82226
rect 347040 82170 361930 82226
rect 361986 82170 362054 82226
rect 362110 82170 362178 82226
rect 362234 82170 362302 82226
rect 362358 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 408594 82226
rect 408650 82170 408718 82226
rect 408774 82170 408842 82226
rect 408898 82170 408966 82226
rect 409022 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 446612 82226
rect 446668 82170 446736 82226
rect 446792 82170 446860 82226
rect 446916 82170 446984 82226
rect 447040 82170 461930 82226
rect 461986 82170 462054 82226
rect 462110 82170 462178 82226
rect 462234 82170 462302 82226
rect 462358 82170 470034 82226
rect 470090 82170 470158 82226
rect 470214 82170 470282 82226
rect 470338 82170 470406 82226
rect 470462 82170 500754 82226
rect 500810 82170 500878 82226
rect 500934 82170 501002 82226
rect 501058 82170 501126 82226
rect 501182 82170 531474 82226
rect 531530 82170 531598 82226
rect 531654 82170 531722 82226
rect 531778 82170 531846 82226
rect 531902 82170 546612 82226
rect 546668 82170 546736 82226
rect 546792 82170 546860 82226
rect 546916 82170 546984 82226
rect 547040 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 61930 82102
rect 61986 82046 62054 82102
rect 62110 82046 62178 82102
rect 62234 82046 62302 82102
rect 62358 82046 70674 82102
rect 70730 82046 70798 82102
rect 70854 82046 70922 82102
rect 70978 82046 71046 82102
rect 71102 82046 101394 82102
rect 101450 82046 101518 82102
rect 101574 82046 101642 82102
rect 101698 82046 101766 82102
rect 101822 82046 132114 82102
rect 132170 82046 132238 82102
rect 132294 82046 132362 82102
rect 132418 82046 132486 82102
rect 132542 82046 146612 82102
rect 146668 82046 146736 82102
rect 146792 82046 146860 82102
rect 146916 82046 146984 82102
rect 147040 82046 161930 82102
rect 161986 82046 162054 82102
rect 162110 82046 162178 82102
rect 162234 82046 162302 82102
rect 162358 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 224274 82102
rect 224330 82046 224398 82102
rect 224454 82046 224522 82102
rect 224578 82046 224646 82102
rect 224702 82046 246612 82102
rect 246668 82046 246736 82102
rect 246792 82046 246860 82102
rect 246916 82046 246984 82102
rect 247040 82046 254994 82102
rect 255050 82046 255118 82102
rect 255174 82046 255242 82102
rect 255298 82046 255366 82102
rect 255422 82046 261930 82102
rect 261986 82046 262054 82102
rect 262110 82046 262178 82102
rect 262234 82046 262302 82102
rect 262358 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 316434 82102
rect 316490 82046 316558 82102
rect 316614 82046 316682 82102
rect 316738 82046 316806 82102
rect 316862 82046 346612 82102
rect 346668 82046 346736 82102
rect 346792 82046 346860 82102
rect 346916 82046 346984 82102
rect 347040 82046 361930 82102
rect 361986 82046 362054 82102
rect 362110 82046 362178 82102
rect 362234 82046 362302 82102
rect 362358 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 408594 82102
rect 408650 82046 408718 82102
rect 408774 82046 408842 82102
rect 408898 82046 408966 82102
rect 409022 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 446612 82102
rect 446668 82046 446736 82102
rect 446792 82046 446860 82102
rect 446916 82046 446984 82102
rect 447040 82046 461930 82102
rect 461986 82046 462054 82102
rect 462110 82046 462178 82102
rect 462234 82046 462302 82102
rect 462358 82046 470034 82102
rect 470090 82046 470158 82102
rect 470214 82046 470282 82102
rect 470338 82046 470406 82102
rect 470462 82046 500754 82102
rect 500810 82046 500878 82102
rect 500934 82046 501002 82102
rect 501058 82046 501126 82102
rect 501182 82046 531474 82102
rect 531530 82046 531598 82102
rect 531654 82046 531722 82102
rect 531778 82046 531846 82102
rect 531902 82046 546612 82102
rect 546668 82046 546736 82102
rect 546792 82046 546860 82102
rect 546916 82046 546984 82102
rect 547040 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 61930 81978
rect 61986 81922 62054 81978
rect 62110 81922 62178 81978
rect 62234 81922 62302 81978
rect 62358 81922 70674 81978
rect 70730 81922 70798 81978
rect 70854 81922 70922 81978
rect 70978 81922 71046 81978
rect 71102 81922 101394 81978
rect 101450 81922 101518 81978
rect 101574 81922 101642 81978
rect 101698 81922 101766 81978
rect 101822 81922 132114 81978
rect 132170 81922 132238 81978
rect 132294 81922 132362 81978
rect 132418 81922 132486 81978
rect 132542 81922 146612 81978
rect 146668 81922 146736 81978
rect 146792 81922 146860 81978
rect 146916 81922 146984 81978
rect 147040 81922 161930 81978
rect 161986 81922 162054 81978
rect 162110 81922 162178 81978
rect 162234 81922 162302 81978
rect 162358 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 224274 81978
rect 224330 81922 224398 81978
rect 224454 81922 224522 81978
rect 224578 81922 224646 81978
rect 224702 81922 246612 81978
rect 246668 81922 246736 81978
rect 246792 81922 246860 81978
rect 246916 81922 246984 81978
rect 247040 81922 254994 81978
rect 255050 81922 255118 81978
rect 255174 81922 255242 81978
rect 255298 81922 255366 81978
rect 255422 81922 261930 81978
rect 261986 81922 262054 81978
rect 262110 81922 262178 81978
rect 262234 81922 262302 81978
rect 262358 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 316434 81978
rect 316490 81922 316558 81978
rect 316614 81922 316682 81978
rect 316738 81922 316806 81978
rect 316862 81922 346612 81978
rect 346668 81922 346736 81978
rect 346792 81922 346860 81978
rect 346916 81922 346984 81978
rect 347040 81922 361930 81978
rect 361986 81922 362054 81978
rect 362110 81922 362178 81978
rect 362234 81922 362302 81978
rect 362358 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 408594 81978
rect 408650 81922 408718 81978
rect 408774 81922 408842 81978
rect 408898 81922 408966 81978
rect 409022 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 446612 81978
rect 446668 81922 446736 81978
rect 446792 81922 446860 81978
rect 446916 81922 446984 81978
rect 447040 81922 461930 81978
rect 461986 81922 462054 81978
rect 462110 81922 462178 81978
rect 462234 81922 462302 81978
rect 462358 81922 470034 81978
rect 470090 81922 470158 81978
rect 470214 81922 470282 81978
rect 470338 81922 470406 81978
rect 470462 81922 500754 81978
rect 500810 81922 500878 81978
rect 500934 81922 501002 81978
rect 501058 81922 501126 81978
rect 501182 81922 531474 81978
rect 531530 81922 531598 81978
rect 531654 81922 531722 81978
rect 531778 81922 531846 81978
rect 531902 81922 546612 81978
rect 546668 81922 546736 81978
rect 546792 81922 546860 81978
rect 546916 81922 546984 81978
rect 547040 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 61130 76350
rect 61186 76294 61254 76350
rect 61310 76294 61378 76350
rect 61434 76294 61502 76350
rect 61558 76294 66954 76350
rect 67010 76294 67078 76350
rect 67134 76294 67202 76350
rect 67258 76294 67326 76350
rect 67382 76294 97674 76350
rect 97730 76294 97798 76350
rect 97854 76294 97922 76350
rect 97978 76294 98046 76350
rect 98102 76294 128394 76350
rect 128450 76294 128518 76350
rect 128574 76294 128642 76350
rect 128698 76294 128766 76350
rect 128822 76294 145812 76350
rect 145868 76294 145936 76350
rect 145992 76294 146060 76350
rect 146116 76294 146184 76350
rect 146240 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 161130 76350
rect 161186 76294 161254 76350
rect 161310 76294 161378 76350
rect 161434 76294 161502 76350
rect 161558 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 245812 76350
rect 245868 76294 245936 76350
rect 245992 76294 246060 76350
rect 246116 76294 246184 76350
rect 246240 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 261130 76350
rect 261186 76294 261254 76350
rect 261310 76294 261378 76350
rect 261434 76294 261502 76350
rect 261558 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 345812 76350
rect 345868 76294 345936 76350
rect 345992 76294 346060 76350
rect 346116 76294 346184 76350
rect 346240 76294 361130 76350
rect 361186 76294 361254 76350
rect 361310 76294 361378 76350
rect 361434 76294 361502 76350
rect 361558 76294 374154 76350
rect 374210 76294 374278 76350
rect 374334 76294 374402 76350
rect 374458 76294 374526 76350
rect 374582 76294 404874 76350
rect 404930 76294 404998 76350
rect 405054 76294 405122 76350
rect 405178 76294 405246 76350
rect 405302 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 445812 76350
rect 445868 76294 445936 76350
rect 445992 76294 446060 76350
rect 446116 76294 446184 76350
rect 446240 76294 461130 76350
rect 461186 76294 461254 76350
rect 461310 76294 461378 76350
rect 461434 76294 461502 76350
rect 461558 76294 466314 76350
rect 466370 76294 466438 76350
rect 466494 76294 466562 76350
rect 466618 76294 466686 76350
rect 466742 76294 497034 76350
rect 497090 76294 497158 76350
rect 497214 76294 497282 76350
rect 497338 76294 497406 76350
rect 497462 76294 527754 76350
rect 527810 76294 527878 76350
rect 527934 76294 528002 76350
rect 528058 76294 528126 76350
rect 528182 76294 545812 76350
rect 545868 76294 545936 76350
rect 545992 76294 546060 76350
rect 546116 76294 546184 76350
rect 546240 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 61130 76226
rect 61186 76170 61254 76226
rect 61310 76170 61378 76226
rect 61434 76170 61502 76226
rect 61558 76170 66954 76226
rect 67010 76170 67078 76226
rect 67134 76170 67202 76226
rect 67258 76170 67326 76226
rect 67382 76170 97674 76226
rect 97730 76170 97798 76226
rect 97854 76170 97922 76226
rect 97978 76170 98046 76226
rect 98102 76170 128394 76226
rect 128450 76170 128518 76226
rect 128574 76170 128642 76226
rect 128698 76170 128766 76226
rect 128822 76170 145812 76226
rect 145868 76170 145936 76226
rect 145992 76170 146060 76226
rect 146116 76170 146184 76226
rect 146240 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 161130 76226
rect 161186 76170 161254 76226
rect 161310 76170 161378 76226
rect 161434 76170 161502 76226
rect 161558 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 245812 76226
rect 245868 76170 245936 76226
rect 245992 76170 246060 76226
rect 246116 76170 246184 76226
rect 246240 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 261130 76226
rect 261186 76170 261254 76226
rect 261310 76170 261378 76226
rect 261434 76170 261502 76226
rect 261558 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 345812 76226
rect 345868 76170 345936 76226
rect 345992 76170 346060 76226
rect 346116 76170 346184 76226
rect 346240 76170 361130 76226
rect 361186 76170 361254 76226
rect 361310 76170 361378 76226
rect 361434 76170 361502 76226
rect 361558 76170 374154 76226
rect 374210 76170 374278 76226
rect 374334 76170 374402 76226
rect 374458 76170 374526 76226
rect 374582 76170 404874 76226
rect 404930 76170 404998 76226
rect 405054 76170 405122 76226
rect 405178 76170 405246 76226
rect 405302 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 445812 76226
rect 445868 76170 445936 76226
rect 445992 76170 446060 76226
rect 446116 76170 446184 76226
rect 446240 76170 461130 76226
rect 461186 76170 461254 76226
rect 461310 76170 461378 76226
rect 461434 76170 461502 76226
rect 461558 76170 466314 76226
rect 466370 76170 466438 76226
rect 466494 76170 466562 76226
rect 466618 76170 466686 76226
rect 466742 76170 497034 76226
rect 497090 76170 497158 76226
rect 497214 76170 497282 76226
rect 497338 76170 497406 76226
rect 497462 76170 527754 76226
rect 527810 76170 527878 76226
rect 527934 76170 528002 76226
rect 528058 76170 528126 76226
rect 528182 76170 545812 76226
rect 545868 76170 545936 76226
rect 545992 76170 546060 76226
rect 546116 76170 546184 76226
rect 546240 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 61130 76102
rect 61186 76046 61254 76102
rect 61310 76046 61378 76102
rect 61434 76046 61502 76102
rect 61558 76046 66954 76102
rect 67010 76046 67078 76102
rect 67134 76046 67202 76102
rect 67258 76046 67326 76102
rect 67382 76046 97674 76102
rect 97730 76046 97798 76102
rect 97854 76046 97922 76102
rect 97978 76046 98046 76102
rect 98102 76046 128394 76102
rect 128450 76046 128518 76102
rect 128574 76046 128642 76102
rect 128698 76046 128766 76102
rect 128822 76046 145812 76102
rect 145868 76046 145936 76102
rect 145992 76046 146060 76102
rect 146116 76046 146184 76102
rect 146240 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 161130 76102
rect 161186 76046 161254 76102
rect 161310 76046 161378 76102
rect 161434 76046 161502 76102
rect 161558 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 245812 76102
rect 245868 76046 245936 76102
rect 245992 76046 246060 76102
rect 246116 76046 246184 76102
rect 246240 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 261130 76102
rect 261186 76046 261254 76102
rect 261310 76046 261378 76102
rect 261434 76046 261502 76102
rect 261558 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 345812 76102
rect 345868 76046 345936 76102
rect 345992 76046 346060 76102
rect 346116 76046 346184 76102
rect 346240 76046 361130 76102
rect 361186 76046 361254 76102
rect 361310 76046 361378 76102
rect 361434 76046 361502 76102
rect 361558 76046 374154 76102
rect 374210 76046 374278 76102
rect 374334 76046 374402 76102
rect 374458 76046 374526 76102
rect 374582 76046 404874 76102
rect 404930 76046 404998 76102
rect 405054 76046 405122 76102
rect 405178 76046 405246 76102
rect 405302 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 445812 76102
rect 445868 76046 445936 76102
rect 445992 76046 446060 76102
rect 446116 76046 446184 76102
rect 446240 76046 461130 76102
rect 461186 76046 461254 76102
rect 461310 76046 461378 76102
rect 461434 76046 461502 76102
rect 461558 76046 466314 76102
rect 466370 76046 466438 76102
rect 466494 76046 466562 76102
rect 466618 76046 466686 76102
rect 466742 76046 497034 76102
rect 497090 76046 497158 76102
rect 497214 76046 497282 76102
rect 497338 76046 497406 76102
rect 497462 76046 527754 76102
rect 527810 76046 527878 76102
rect 527934 76046 528002 76102
rect 528058 76046 528126 76102
rect 528182 76046 545812 76102
rect 545868 76046 545936 76102
rect 545992 76046 546060 76102
rect 546116 76046 546184 76102
rect 546240 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 61130 75978
rect 61186 75922 61254 75978
rect 61310 75922 61378 75978
rect 61434 75922 61502 75978
rect 61558 75922 66954 75978
rect 67010 75922 67078 75978
rect 67134 75922 67202 75978
rect 67258 75922 67326 75978
rect 67382 75922 97674 75978
rect 97730 75922 97798 75978
rect 97854 75922 97922 75978
rect 97978 75922 98046 75978
rect 98102 75922 128394 75978
rect 128450 75922 128518 75978
rect 128574 75922 128642 75978
rect 128698 75922 128766 75978
rect 128822 75922 145812 75978
rect 145868 75922 145936 75978
rect 145992 75922 146060 75978
rect 146116 75922 146184 75978
rect 146240 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 161130 75978
rect 161186 75922 161254 75978
rect 161310 75922 161378 75978
rect 161434 75922 161502 75978
rect 161558 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 245812 75978
rect 245868 75922 245936 75978
rect 245992 75922 246060 75978
rect 246116 75922 246184 75978
rect 246240 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 261130 75978
rect 261186 75922 261254 75978
rect 261310 75922 261378 75978
rect 261434 75922 261502 75978
rect 261558 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 345812 75978
rect 345868 75922 345936 75978
rect 345992 75922 346060 75978
rect 346116 75922 346184 75978
rect 346240 75922 361130 75978
rect 361186 75922 361254 75978
rect 361310 75922 361378 75978
rect 361434 75922 361502 75978
rect 361558 75922 374154 75978
rect 374210 75922 374278 75978
rect 374334 75922 374402 75978
rect 374458 75922 374526 75978
rect 374582 75922 404874 75978
rect 404930 75922 404998 75978
rect 405054 75922 405122 75978
rect 405178 75922 405246 75978
rect 405302 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 445812 75978
rect 445868 75922 445936 75978
rect 445992 75922 446060 75978
rect 446116 75922 446184 75978
rect 446240 75922 461130 75978
rect 461186 75922 461254 75978
rect 461310 75922 461378 75978
rect 461434 75922 461502 75978
rect 461558 75922 466314 75978
rect 466370 75922 466438 75978
rect 466494 75922 466562 75978
rect 466618 75922 466686 75978
rect 466742 75922 497034 75978
rect 497090 75922 497158 75978
rect 497214 75922 497282 75978
rect 497338 75922 497406 75978
rect 497462 75922 527754 75978
rect 527810 75922 527878 75978
rect 527934 75922 528002 75978
rect 528058 75922 528126 75978
rect 528182 75922 545812 75978
rect 545868 75922 545936 75978
rect 545992 75922 546060 75978
rect 546116 75922 546184 75978
rect 546240 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 61930 64350
rect 61986 64294 62054 64350
rect 62110 64294 62178 64350
rect 62234 64294 62302 64350
rect 62358 64294 70674 64350
rect 70730 64294 70798 64350
rect 70854 64294 70922 64350
rect 70978 64294 71046 64350
rect 71102 64294 101394 64350
rect 101450 64294 101518 64350
rect 101574 64294 101642 64350
rect 101698 64294 101766 64350
rect 101822 64294 132114 64350
rect 132170 64294 132238 64350
rect 132294 64294 132362 64350
rect 132418 64294 132486 64350
rect 132542 64294 146612 64350
rect 146668 64294 146736 64350
rect 146792 64294 146860 64350
rect 146916 64294 146984 64350
rect 147040 64294 161930 64350
rect 161986 64294 162054 64350
rect 162110 64294 162178 64350
rect 162234 64294 162302 64350
rect 162358 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 193554 64350
rect 193610 64294 193678 64350
rect 193734 64294 193802 64350
rect 193858 64294 193926 64350
rect 193982 64294 224274 64350
rect 224330 64294 224398 64350
rect 224454 64294 224522 64350
rect 224578 64294 224646 64350
rect 224702 64294 246612 64350
rect 246668 64294 246736 64350
rect 246792 64294 246860 64350
rect 246916 64294 246984 64350
rect 247040 64294 254994 64350
rect 255050 64294 255118 64350
rect 255174 64294 255242 64350
rect 255298 64294 255366 64350
rect 255422 64294 261930 64350
rect 261986 64294 262054 64350
rect 262110 64294 262178 64350
rect 262234 64294 262302 64350
rect 262358 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 316434 64350
rect 316490 64294 316558 64350
rect 316614 64294 316682 64350
rect 316738 64294 316806 64350
rect 316862 64294 346612 64350
rect 346668 64294 346736 64350
rect 346792 64294 346860 64350
rect 346916 64294 346984 64350
rect 347040 64294 361930 64350
rect 361986 64294 362054 64350
rect 362110 64294 362178 64350
rect 362234 64294 362302 64350
rect 362358 64294 377874 64350
rect 377930 64294 377998 64350
rect 378054 64294 378122 64350
rect 378178 64294 378246 64350
rect 378302 64294 408594 64350
rect 408650 64294 408718 64350
rect 408774 64294 408842 64350
rect 408898 64294 408966 64350
rect 409022 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 446612 64350
rect 446668 64294 446736 64350
rect 446792 64294 446860 64350
rect 446916 64294 446984 64350
rect 447040 64294 461930 64350
rect 461986 64294 462054 64350
rect 462110 64294 462178 64350
rect 462234 64294 462302 64350
rect 462358 64294 470034 64350
rect 470090 64294 470158 64350
rect 470214 64294 470282 64350
rect 470338 64294 470406 64350
rect 470462 64294 500754 64350
rect 500810 64294 500878 64350
rect 500934 64294 501002 64350
rect 501058 64294 501126 64350
rect 501182 64294 531474 64350
rect 531530 64294 531598 64350
rect 531654 64294 531722 64350
rect 531778 64294 531846 64350
rect 531902 64294 546612 64350
rect 546668 64294 546736 64350
rect 546792 64294 546860 64350
rect 546916 64294 546984 64350
rect 547040 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 61930 64226
rect 61986 64170 62054 64226
rect 62110 64170 62178 64226
rect 62234 64170 62302 64226
rect 62358 64170 70674 64226
rect 70730 64170 70798 64226
rect 70854 64170 70922 64226
rect 70978 64170 71046 64226
rect 71102 64170 101394 64226
rect 101450 64170 101518 64226
rect 101574 64170 101642 64226
rect 101698 64170 101766 64226
rect 101822 64170 132114 64226
rect 132170 64170 132238 64226
rect 132294 64170 132362 64226
rect 132418 64170 132486 64226
rect 132542 64170 146612 64226
rect 146668 64170 146736 64226
rect 146792 64170 146860 64226
rect 146916 64170 146984 64226
rect 147040 64170 161930 64226
rect 161986 64170 162054 64226
rect 162110 64170 162178 64226
rect 162234 64170 162302 64226
rect 162358 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 193554 64226
rect 193610 64170 193678 64226
rect 193734 64170 193802 64226
rect 193858 64170 193926 64226
rect 193982 64170 224274 64226
rect 224330 64170 224398 64226
rect 224454 64170 224522 64226
rect 224578 64170 224646 64226
rect 224702 64170 246612 64226
rect 246668 64170 246736 64226
rect 246792 64170 246860 64226
rect 246916 64170 246984 64226
rect 247040 64170 254994 64226
rect 255050 64170 255118 64226
rect 255174 64170 255242 64226
rect 255298 64170 255366 64226
rect 255422 64170 261930 64226
rect 261986 64170 262054 64226
rect 262110 64170 262178 64226
rect 262234 64170 262302 64226
rect 262358 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 316434 64226
rect 316490 64170 316558 64226
rect 316614 64170 316682 64226
rect 316738 64170 316806 64226
rect 316862 64170 346612 64226
rect 346668 64170 346736 64226
rect 346792 64170 346860 64226
rect 346916 64170 346984 64226
rect 347040 64170 361930 64226
rect 361986 64170 362054 64226
rect 362110 64170 362178 64226
rect 362234 64170 362302 64226
rect 362358 64170 377874 64226
rect 377930 64170 377998 64226
rect 378054 64170 378122 64226
rect 378178 64170 378246 64226
rect 378302 64170 408594 64226
rect 408650 64170 408718 64226
rect 408774 64170 408842 64226
rect 408898 64170 408966 64226
rect 409022 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 446612 64226
rect 446668 64170 446736 64226
rect 446792 64170 446860 64226
rect 446916 64170 446984 64226
rect 447040 64170 461930 64226
rect 461986 64170 462054 64226
rect 462110 64170 462178 64226
rect 462234 64170 462302 64226
rect 462358 64170 470034 64226
rect 470090 64170 470158 64226
rect 470214 64170 470282 64226
rect 470338 64170 470406 64226
rect 470462 64170 500754 64226
rect 500810 64170 500878 64226
rect 500934 64170 501002 64226
rect 501058 64170 501126 64226
rect 501182 64170 531474 64226
rect 531530 64170 531598 64226
rect 531654 64170 531722 64226
rect 531778 64170 531846 64226
rect 531902 64170 546612 64226
rect 546668 64170 546736 64226
rect 546792 64170 546860 64226
rect 546916 64170 546984 64226
rect 547040 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 61930 64102
rect 61986 64046 62054 64102
rect 62110 64046 62178 64102
rect 62234 64046 62302 64102
rect 62358 64046 70674 64102
rect 70730 64046 70798 64102
rect 70854 64046 70922 64102
rect 70978 64046 71046 64102
rect 71102 64046 101394 64102
rect 101450 64046 101518 64102
rect 101574 64046 101642 64102
rect 101698 64046 101766 64102
rect 101822 64046 132114 64102
rect 132170 64046 132238 64102
rect 132294 64046 132362 64102
rect 132418 64046 132486 64102
rect 132542 64046 146612 64102
rect 146668 64046 146736 64102
rect 146792 64046 146860 64102
rect 146916 64046 146984 64102
rect 147040 64046 161930 64102
rect 161986 64046 162054 64102
rect 162110 64046 162178 64102
rect 162234 64046 162302 64102
rect 162358 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 193554 64102
rect 193610 64046 193678 64102
rect 193734 64046 193802 64102
rect 193858 64046 193926 64102
rect 193982 64046 224274 64102
rect 224330 64046 224398 64102
rect 224454 64046 224522 64102
rect 224578 64046 224646 64102
rect 224702 64046 246612 64102
rect 246668 64046 246736 64102
rect 246792 64046 246860 64102
rect 246916 64046 246984 64102
rect 247040 64046 254994 64102
rect 255050 64046 255118 64102
rect 255174 64046 255242 64102
rect 255298 64046 255366 64102
rect 255422 64046 261930 64102
rect 261986 64046 262054 64102
rect 262110 64046 262178 64102
rect 262234 64046 262302 64102
rect 262358 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 316434 64102
rect 316490 64046 316558 64102
rect 316614 64046 316682 64102
rect 316738 64046 316806 64102
rect 316862 64046 346612 64102
rect 346668 64046 346736 64102
rect 346792 64046 346860 64102
rect 346916 64046 346984 64102
rect 347040 64046 361930 64102
rect 361986 64046 362054 64102
rect 362110 64046 362178 64102
rect 362234 64046 362302 64102
rect 362358 64046 377874 64102
rect 377930 64046 377998 64102
rect 378054 64046 378122 64102
rect 378178 64046 378246 64102
rect 378302 64046 408594 64102
rect 408650 64046 408718 64102
rect 408774 64046 408842 64102
rect 408898 64046 408966 64102
rect 409022 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 446612 64102
rect 446668 64046 446736 64102
rect 446792 64046 446860 64102
rect 446916 64046 446984 64102
rect 447040 64046 461930 64102
rect 461986 64046 462054 64102
rect 462110 64046 462178 64102
rect 462234 64046 462302 64102
rect 462358 64046 470034 64102
rect 470090 64046 470158 64102
rect 470214 64046 470282 64102
rect 470338 64046 470406 64102
rect 470462 64046 500754 64102
rect 500810 64046 500878 64102
rect 500934 64046 501002 64102
rect 501058 64046 501126 64102
rect 501182 64046 531474 64102
rect 531530 64046 531598 64102
rect 531654 64046 531722 64102
rect 531778 64046 531846 64102
rect 531902 64046 546612 64102
rect 546668 64046 546736 64102
rect 546792 64046 546860 64102
rect 546916 64046 546984 64102
rect 547040 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 61930 63978
rect 61986 63922 62054 63978
rect 62110 63922 62178 63978
rect 62234 63922 62302 63978
rect 62358 63922 70674 63978
rect 70730 63922 70798 63978
rect 70854 63922 70922 63978
rect 70978 63922 71046 63978
rect 71102 63922 101394 63978
rect 101450 63922 101518 63978
rect 101574 63922 101642 63978
rect 101698 63922 101766 63978
rect 101822 63922 132114 63978
rect 132170 63922 132238 63978
rect 132294 63922 132362 63978
rect 132418 63922 132486 63978
rect 132542 63922 146612 63978
rect 146668 63922 146736 63978
rect 146792 63922 146860 63978
rect 146916 63922 146984 63978
rect 147040 63922 161930 63978
rect 161986 63922 162054 63978
rect 162110 63922 162178 63978
rect 162234 63922 162302 63978
rect 162358 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 193554 63978
rect 193610 63922 193678 63978
rect 193734 63922 193802 63978
rect 193858 63922 193926 63978
rect 193982 63922 224274 63978
rect 224330 63922 224398 63978
rect 224454 63922 224522 63978
rect 224578 63922 224646 63978
rect 224702 63922 246612 63978
rect 246668 63922 246736 63978
rect 246792 63922 246860 63978
rect 246916 63922 246984 63978
rect 247040 63922 254994 63978
rect 255050 63922 255118 63978
rect 255174 63922 255242 63978
rect 255298 63922 255366 63978
rect 255422 63922 261930 63978
rect 261986 63922 262054 63978
rect 262110 63922 262178 63978
rect 262234 63922 262302 63978
rect 262358 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 316434 63978
rect 316490 63922 316558 63978
rect 316614 63922 316682 63978
rect 316738 63922 316806 63978
rect 316862 63922 346612 63978
rect 346668 63922 346736 63978
rect 346792 63922 346860 63978
rect 346916 63922 346984 63978
rect 347040 63922 361930 63978
rect 361986 63922 362054 63978
rect 362110 63922 362178 63978
rect 362234 63922 362302 63978
rect 362358 63922 377874 63978
rect 377930 63922 377998 63978
rect 378054 63922 378122 63978
rect 378178 63922 378246 63978
rect 378302 63922 408594 63978
rect 408650 63922 408718 63978
rect 408774 63922 408842 63978
rect 408898 63922 408966 63978
rect 409022 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 446612 63978
rect 446668 63922 446736 63978
rect 446792 63922 446860 63978
rect 446916 63922 446984 63978
rect 447040 63922 461930 63978
rect 461986 63922 462054 63978
rect 462110 63922 462178 63978
rect 462234 63922 462302 63978
rect 462358 63922 470034 63978
rect 470090 63922 470158 63978
rect 470214 63922 470282 63978
rect 470338 63922 470406 63978
rect 470462 63922 500754 63978
rect 500810 63922 500878 63978
rect 500934 63922 501002 63978
rect 501058 63922 501126 63978
rect 501182 63922 531474 63978
rect 531530 63922 531598 63978
rect 531654 63922 531722 63978
rect 531778 63922 531846 63978
rect 531902 63922 546612 63978
rect 546668 63922 546736 63978
rect 546792 63922 546860 63978
rect 546916 63922 546984 63978
rect 547040 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 61130 58350
rect 61186 58294 61254 58350
rect 61310 58294 61378 58350
rect 61434 58294 61502 58350
rect 61558 58294 66954 58350
rect 67010 58294 67078 58350
rect 67134 58294 67202 58350
rect 67258 58294 67326 58350
rect 67382 58294 97674 58350
rect 97730 58294 97798 58350
rect 97854 58294 97922 58350
rect 97978 58294 98046 58350
rect 98102 58294 128394 58350
rect 128450 58294 128518 58350
rect 128574 58294 128642 58350
rect 128698 58294 128766 58350
rect 128822 58294 145812 58350
rect 145868 58294 145936 58350
rect 145992 58294 146060 58350
rect 146116 58294 146184 58350
rect 146240 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 161130 58350
rect 161186 58294 161254 58350
rect 161310 58294 161378 58350
rect 161434 58294 161502 58350
rect 161558 58294 189834 58350
rect 189890 58294 189958 58350
rect 190014 58294 190082 58350
rect 190138 58294 190206 58350
rect 190262 58294 220554 58350
rect 220610 58294 220678 58350
rect 220734 58294 220802 58350
rect 220858 58294 220926 58350
rect 220982 58294 245812 58350
rect 245868 58294 245936 58350
rect 245992 58294 246060 58350
rect 246116 58294 246184 58350
rect 246240 58294 251274 58350
rect 251330 58294 251398 58350
rect 251454 58294 251522 58350
rect 251578 58294 251646 58350
rect 251702 58294 261130 58350
rect 261186 58294 261254 58350
rect 261310 58294 261378 58350
rect 261434 58294 261502 58350
rect 261558 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 345812 58350
rect 345868 58294 345936 58350
rect 345992 58294 346060 58350
rect 346116 58294 346184 58350
rect 346240 58294 361130 58350
rect 361186 58294 361254 58350
rect 361310 58294 361378 58350
rect 361434 58294 361502 58350
rect 361558 58294 374154 58350
rect 374210 58294 374278 58350
rect 374334 58294 374402 58350
rect 374458 58294 374526 58350
rect 374582 58294 404874 58350
rect 404930 58294 404998 58350
rect 405054 58294 405122 58350
rect 405178 58294 405246 58350
rect 405302 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 445812 58350
rect 445868 58294 445936 58350
rect 445992 58294 446060 58350
rect 446116 58294 446184 58350
rect 446240 58294 461130 58350
rect 461186 58294 461254 58350
rect 461310 58294 461378 58350
rect 461434 58294 461502 58350
rect 461558 58294 466314 58350
rect 466370 58294 466438 58350
rect 466494 58294 466562 58350
rect 466618 58294 466686 58350
rect 466742 58294 497034 58350
rect 497090 58294 497158 58350
rect 497214 58294 497282 58350
rect 497338 58294 497406 58350
rect 497462 58294 527754 58350
rect 527810 58294 527878 58350
rect 527934 58294 528002 58350
rect 528058 58294 528126 58350
rect 528182 58294 545812 58350
rect 545868 58294 545936 58350
rect 545992 58294 546060 58350
rect 546116 58294 546184 58350
rect 546240 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 61130 58226
rect 61186 58170 61254 58226
rect 61310 58170 61378 58226
rect 61434 58170 61502 58226
rect 61558 58170 66954 58226
rect 67010 58170 67078 58226
rect 67134 58170 67202 58226
rect 67258 58170 67326 58226
rect 67382 58170 97674 58226
rect 97730 58170 97798 58226
rect 97854 58170 97922 58226
rect 97978 58170 98046 58226
rect 98102 58170 128394 58226
rect 128450 58170 128518 58226
rect 128574 58170 128642 58226
rect 128698 58170 128766 58226
rect 128822 58170 145812 58226
rect 145868 58170 145936 58226
rect 145992 58170 146060 58226
rect 146116 58170 146184 58226
rect 146240 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 161130 58226
rect 161186 58170 161254 58226
rect 161310 58170 161378 58226
rect 161434 58170 161502 58226
rect 161558 58170 189834 58226
rect 189890 58170 189958 58226
rect 190014 58170 190082 58226
rect 190138 58170 190206 58226
rect 190262 58170 220554 58226
rect 220610 58170 220678 58226
rect 220734 58170 220802 58226
rect 220858 58170 220926 58226
rect 220982 58170 245812 58226
rect 245868 58170 245936 58226
rect 245992 58170 246060 58226
rect 246116 58170 246184 58226
rect 246240 58170 251274 58226
rect 251330 58170 251398 58226
rect 251454 58170 251522 58226
rect 251578 58170 251646 58226
rect 251702 58170 261130 58226
rect 261186 58170 261254 58226
rect 261310 58170 261378 58226
rect 261434 58170 261502 58226
rect 261558 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 345812 58226
rect 345868 58170 345936 58226
rect 345992 58170 346060 58226
rect 346116 58170 346184 58226
rect 346240 58170 361130 58226
rect 361186 58170 361254 58226
rect 361310 58170 361378 58226
rect 361434 58170 361502 58226
rect 361558 58170 374154 58226
rect 374210 58170 374278 58226
rect 374334 58170 374402 58226
rect 374458 58170 374526 58226
rect 374582 58170 404874 58226
rect 404930 58170 404998 58226
rect 405054 58170 405122 58226
rect 405178 58170 405246 58226
rect 405302 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 445812 58226
rect 445868 58170 445936 58226
rect 445992 58170 446060 58226
rect 446116 58170 446184 58226
rect 446240 58170 461130 58226
rect 461186 58170 461254 58226
rect 461310 58170 461378 58226
rect 461434 58170 461502 58226
rect 461558 58170 466314 58226
rect 466370 58170 466438 58226
rect 466494 58170 466562 58226
rect 466618 58170 466686 58226
rect 466742 58170 497034 58226
rect 497090 58170 497158 58226
rect 497214 58170 497282 58226
rect 497338 58170 497406 58226
rect 497462 58170 527754 58226
rect 527810 58170 527878 58226
rect 527934 58170 528002 58226
rect 528058 58170 528126 58226
rect 528182 58170 545812 58226
rect 545868 58170 545936 58226
rect 545992 58170 546060 58226
rect 546116 58170 546184 58226
rect 546240 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 61130 58102
rect 61186 58046 61254 58102
rect 61310 58046 61378 58102
rect 61434 58046 61502 58102
rect 61558 58046 66954 58102
rect 67010 58046 67078 58102
rect 67134 58046 67202 58102
rect 67258 58046 67326 58102
rect 67382 58046 97674 58102
rect 97730 58046 97798 58102
rect 97854 58046 97922 58102
rect 97978 58046 98046 58102
rect 98102 58046 128394 58102
rect 128450 58046 128518 58102
rect 128574 58046 128642 58102
rect 128698 58046 128766 58102
rect 128822 58046 145812 58102
rect 145868 58046 145936 58102
rect 145992 58046 146060 58102
rect 146116 58046 146184 58102
rect 146240 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 161130 58102
rect 161186 58046 161254 58102
rect 161310 58046 161378 58102
rect 161434 58046 161502 58102
rect 161558 58046 189834 58102
rect 189890 58046 189958 58102
rect 190014 58046 190082 58102
rect 190138 58046 190206 58102
rect 190262 58046 220554 58102
rect 220610 58046 220678 58102
rect 220734 58046 220802 58102
rect 220858 58046 220926 58102
rect 220982 58046 245812 58102
rect 245868 58046 245936 58102
rect 245992 58046 246060 58102
rect 246116 58046 246184 58102
rect 246240 58046 251274 58102
rect 251330 58046 251398 58102
rect 251454 58046 251522 58102
rect 251578 58046 251646 58102
rect 251702 58046 261130 58102
rect 261186 58046 261254 58102
rect 261310 58046 261378 58102
rect 261434 58046 261502 58102
rect 261558 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 345812 58102
rect 345868 58046 345936 58102
rect 345992 58046 346060 58102
rect 346116 58046 346184 58102
rect 346240 58046 361130 58102
rect 361186 58046 361254 58102
rect 361310 58046 361378 58102
rect 361434 58046 361502 58102
rect 361558 58046 374154 58102
rect 374210 58046 374278 58102
rect 374334 58046 374402 58102
rect 374458 58046 374526 58102
rect 374582 58046 404874 58102
rect 404930 58046 404998 58102
rect 405054 58046 405122 58102
rect 405178 58046 405246 58102
rect 405302 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 445812 58102
rect 445868 58046 445936 58102
rect 445992 58046 446060 58102
rect 446116 58046 446184 58102
rect 446240 58046 461130 58102
rect 461186 58046 461254 58102
rect 461310 58046 461378 58102
rect 461434 58046 461502 58102
rect 461558 58046 466314 58102
rect 466370 58046 466438 58102
rect 466494 58046 466562 58102
rect 466618 58046 466686 58102
rect 466742 58046 497034 58102
rect 497090 58046 497158 58102
rect 497214 58046 497282 58102
rect 497338 58046 497406 58102
rect 497462 58046 527754 58102
rect 527810 58046 527878 58102
rect 527934 58046 528002 58102
rect 528058 58046 528126 58102
rect 528182 58046 545812 58102
rect 545868 58046 545936 58102
rect 545992 58046 546060 58102
rect 546116 58046 546184 58102
rect 546240 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 61130 57978
rect 61186 57922 61254 57978
rect 61310 57922 61378 57978
rect 61434 57922 61502 57978
rect 61558 57922 66954 57978
rect 67010 57922 67078 57978
rect 67134 57922 67202 57978
rect 67258 57922 67326 57978
rect 67382 57922 97674 57978
rect 97730 57922 97798 57978
rect 97854 57922 97922 57978
rect 97978 57922 98046 57978
rect 98102 57922 128394 57978
rect 128450 57922 128518 57978
rect 128574 57922 128642 57978
rect 128698 57922 128766 57978
rect 128822 57922 145812 57978
rect 145868 57922 145936 57978
rect 145992 57922 146060 57978
rect 146116 57922 146184 57978
rect 146240 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 161130 57978
rect 161186 57922 161254 57978
rect 161310 57922 161378 57978
rect 161434 57922 161502 57978
rect 161558 57922 189834 57978
rect 189890 57922 189958 57978
rect 190014 57922 190082 57978
rect 190138 57922 190206 57978
rect 190262 57922 220554 57978
rect 220610 57922 220678 57978
rect 220734 57922 220802 57978
rect 220858 57922 220926 57978
rect 220982 57922 245812 57978
rect 245868 57922 245936 57978
rect 245992 57922 246060 57978
rect 246116 57922 246184 57978
rect 246240 57922 251274 57978
rect 251330 57922 251398 57978
rect 251454 57922 251522 57978
rect 251578 57922 251646 57978
rect 251702 57922 261130 57978
rect 261186 57922 261254 57978
rect 261310 57922 261378 57978
rect 261434 57922 261502 57978
rect 261558 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 345812 57978
rect 345868 57922 345936 57978
rect 345992 57922 346060 57978
rect 346116 57922 346184 57978
rect 346240 57922 361130 57978
rect 361186 57922 361254 57978
rect 361310 57922 361378 57978
rect 361434 57922 361502 57978
rect 361558 57922 374154 57978
rect 374210 57922 374278 57978
rect 374334 57922 374402 57978
rect 374458 57922 374526 57978
rect 374582 57922 404874 57978
rect 404930 57922 404998 57978
rect 405054 57922 405122 57978
rect 405178 57922 405246 57978
rect 405302 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 445812 57978
rect 445868 57922 445936 57978
rect 445992 57922 446060 57978
rect 446116 57922 446184 57978
rect 446240 57922 461130 57978
rect 461186 57922 461254 57978
rect 461310 57922 461378 57978
rect 461434 57922 461502 57978
rect 461558 57922 466314 57978
rect 466370 57922 466438 57978
rect 466494 57922 466562 57978
rect 466618 57922 466686 57978
rect 466742 57922 497034 57978
rect 497090 57922 497158 57978
rect 497214 57922 497282 57978
rect 497338 57922 497406 57978
rect 497462 57922 527754 57978
rect 527810 57922 527878 57978
rect 527934 57922 528002 57978
rect 528058 57922 528126 57978
rect 528182 57922 545812 57978
rect 545868 57922 545936 57978
rect 545992 57922 546060 57978
rect 546116 57922 546184 57978
rect 546240 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 61930 46350
rect 61986 46294 62054 46350
rect 62110 46294 62178 46350
rect 62234 46294 62302 46350
rect 62358 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 146612 46350
rect 146668 46294 146736 46350
rect 146792 46294 146860 46350
rect 146916 46294 146984 46350
rect 147040 46294 161930 46350
rect 161986 46294 162054 46350
rect 162110 46294 162178 46350
rect 162234 46294 162302 46350
rect 162358 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 246612 46350
rect 246668 46294 246736 46350
rect 246792 46294 246860 46350
rect 246916 46294 246984 46350
rect 247040 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 261930 46350
rect 261986 46294 262054 46350
rect 262110 46294 262178 46350
rect 262234 46294 262302 46350
rect 262358 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 346612 46350
rect 346668 46294 346736 46350
rect 346792 46294 346860 46350
rect 346916 46294 346984 46350
rect 347040 46294 361930 46350
rect 361986 46294 362054 46350
rect 362110 46294 362178 46350
rect 362234 46294 362302 46350
rect 362358 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 446612 46350
rect 446668 46294 446736 46350
rect 446792 46294 446860 46350
rect 446916 46294 446984 46350
rect 447040 46294 461930 46350
rect 461986 46294 462054 46350
rect 462110 46294 462178 46350
rect 462234 46294 462302 46350
rect 462358 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 546612 46350
rect 546668 46294 546736 46350
rect 546792 46294 546860 46350
rect 546916 46294 546984 46350
rect 547040 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 61930 46226
rect 61986 46170 62054 46226
rect 62110 46170 62178 46226
rect 62234 46170 62302 46226
rect 62358 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 146612 46226
rect 146668 46170 146736 46226
rect 146792 46170 146860 46226
rect 146916 46170 146984 46226
rect 147040 46170 161930 46226
rect 161986 46170 162054 46226
rect 162110 46170 162178 46226
rect 162234 46170 162302 46226
rect 162358 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 246612 46226
rect 246668 46170 246736 46226
rect 246792 46170 246860 46226
rect 246916 46170 246984 46226
rect 247040 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 261930 46226
rect 261986 46170 262054 46226
rect 262110 46170 262178 46226
rect 262234 46170 262302 46226
rect 262358 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 346612 46226
rect 346668 46170 346736 46226
rect 346792 46170 346860 46226
rect 346916 46170 346984 46226
rect 347040 46170 361930 46226
rect 361986 46170 362054 46226
rect 362110 46170 362178 46226
rect 362234 46170 362302 46226
rect 362358 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 446612 46226
rect 446668 46170 446736 46226
rect 446792 46170 446860 46226
rect 446916 46170 446984 46226
rect 447040 46170 461930 46226
rect 461986 46170 462054 46226
rect 462110 46170 462178 46226
rect 462234 46170 462302 46226
rect 462358 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 546612 46226
rect 546668 46170 546736 46226
rect 546792 46170 546860 46226
rect 546916 46170 546984 46226
rect 547040 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 61930 46102
rect 61986 46046 62054 46102
rect 62110 46046 62178 46102
rect 62234 46046 62302 46102
rect 62358 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 146612 46102
rect 146668 46046 146736 46102
rect 146792 46046 146860 46102
rect 146916 46046 146984 46102
rect 147040 46046 161930 46102
rect 161986 46046 162054 46102
rect 162110 46046 162178 46102
rect 162234 46046 162302 46102
rect 162358 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 246612 46102
rect 246668 46046 246736 46102
rect 246792 46046 246860 46102
rect 246916 46046 246984 46102
rect 247040 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 261930 46102
rect 261986 46046 262054 46102
rect 262110 46046 262178 46102
rect 262234 46046 262302 46102
rect 262358 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 346612 46102
rect 346668 46046 346736 46102
rect 346792 46046 346860 46102
rect 346916 46046 346984 46102
rect 347040 46046 361930 46102
rect 361986 46046 362054 46102
rect 362110 46046 362178 46102
rect 362234 46046 362302 46102
rect 362358 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 446612 46102
rect 446668 46046 446736 46102
rect 446792 46046 446860 46102
rect 446916 46046 446984 46102
rect 447040 46046 461930 46102
rect 461986 46046 462054 46102
rect 462110 46046 462178 46102
rect 462234 46046 462302 46102
rect 462358 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 546612 46102
rect 546668 46046 546736 46102
rect 546792 46046 546860 46102
rect 546916 46046 546984 46102
rect 547040 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 61930 45978
rect 61986 45922 62054 45978
rect 62110 45922 62178 45978
rect 62234 45922 62302 45978
rect 62358 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 146612 45978
rect 146668 45922 146736 45978
rect 146792 45922 146860 45978
rect 146916 45922 146984 45978
rect 147040 45922 161930 45978
rect 161986 45922 162054 45978
rect 162110 45922 162178 45978
rect 162234 45922 162302 45978
rect 162358 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 246612 45978
rect 246668 45922 246736 45978
rect 246792 45922 246860 45978
rect 246916 45922 246984 45978
rect 247040 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 261930 45978
rect 261986 45922 262054 45978
rect 262110 45922 262178 45978
rect 262234 45922 262302 45978
rect 262358 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 346612 45978
rect 346668 45922 346736 45978
rect 346792 45922 346860 45978
rect 346916 45922 346984 45978
rect 347040 45922 361930 45978
rect 361986 45922 362054 45978
rect 362110 45922 362178 45978
rect 362234 45922 362302 45978
rect 362358 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 446612 45978
rect 446668 45922 446736 45978
rect 446792 45922 446860 45978
rect 446916 45922 446984 45978
rect 447040 45922 461930 45978
rect 461986 45922 462054 45978
rect 462110 45922 462178 45978
rect 462234 45922 462302 45978
rect 462358 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 546612 45978
rect 546668 45922 546736 45978
rect 546792 45922 546860 45978
rect 546916 45922 546984 45978
rect 547040 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect 137212 4978 155556 4994
rect 137212 4922 137228 4978
rect 137284 4922 155484 4978
rect 155540 4922 155556 4978
rect 137212 4906 155556 4922
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use avali_logo  avali_logo
timestamp 0
transform 1 0 60000 0 1 490000
box 0 0 60000 70440
use boot_rom  boot_rom
timestamp 0
transform 1 0 480000 0 1 300000
box 0 3076 40656 42000
use gpios  gpios
timestamp 0
transform 1 0 480000 0 1 380000
box 0 0 50000 50000
use ram_controller  ram_controller
timestamp 0
transform 1 0 60000 0 1 160000
box 1258 0 218710 50000
use serial_ports  serial_ports
timestamp 0
transform 1 0 160000 0 1 500000
box 1258 0 55000 55000
use sid_top  sid
timestamp 0
transform 1 0 300000 0 1 400000
box 1250 3076 148624 150000
use gf180_ram_512x8_wrapper_as2650  sram0
timestamp 0
transform 1 0 60000 0 1 40000
box 1000 1000 87372 99176
use gf180_ram_512x8_wrapper_as2650  sram1
timestamp 0
transform 1 0 160000 0 1 40000
box 1000 1000 87372 99176
use gf180_ram_512x8_wrapper_as2650  sram2
timestamp 0
transform 1 0 260000 0 1 40000
box 1000 1000 87372 99176
use gf180_ram_512x8_wrapper_as2650  sram3
timestamp 0
transform 1 0 360000 0 1 40000
box 1000 1000 87372 99176
use gf180_ram_512x8_wrapper_as2650  sram4
timestamp 0
transform 1 0 460000 0 1 40000
box 1000 1000 87372 99176
use gf180_ram_512x8_wrapper_as2650  sram5
timestamp 0
transform -1 0 558972 0 -1 259176
box 1000 1000 87372 99176
use gf180_ram_512x8_wrapper_as2650  sram6
timestamp 0
transform 1 0 360000 0 1 160000
box 1000 1000 87372 99176
use gf180_ram_512x8_wrapper_as2650  sram7
timestamp 0
transform -1 0 388972 0 -1 379176
box 1000 1000 87372 99176
use timers  timers
timestamp 0
transform 1 0 470000 0 1 450000
box 0 0 85000 85000
use wrapped_as2650  wrapped_as2650
timestamp 0
transform 1 0 60000 0 1 290000
box 0 0 210000 140000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 494488 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 533992 67478 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 299890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 425262 98198 490648 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 551392 98198 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 299890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 425262 128918 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 299890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 425262 159638 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 299890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 425262 190358 501266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 548798 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 162274 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 169150 221078 299890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 425262 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 299890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 425262 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 402722 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 548142 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 402722 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 548142 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 402722 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 548142 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 402722 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 548142 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 402722 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 548142 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 305970 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 340062 497558 387426 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 526238 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 453058 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 526238 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 491608 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 536872 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 299890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 425262 101918 493168 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 556192 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 299890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 425262 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 299890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 425262 163358 501266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 548798 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 299890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 425262 194078 501266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 548798 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 162274 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 169150 224798 299890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 425262 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 299890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 425262 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 -1644 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 -1644 316958 402722 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 548142 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 -1644 347678 41024 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 137760 347678 402722 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 548142 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 -1644 378398 402722 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 548142 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 -1644 409118 402722 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 548142 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 402722 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 548142 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 305970 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 340062 501278 387426 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 526238 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 453058 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 526238 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 251674 292322 251674 292322 0 vdd
rlabel via4 264350 424322 264350 424322 0 vss
rlabel metal2 212968 140742 212968 140742 0 A_all\[0\]
rlabel metal2 114744 140126 114744 140126 0 A_all\[1\]
rlabel metal2 116606 139048 116606 139048 0 A_all\[2\]
rlabel metal2 96488 141008 96488 141008 0 A_all\[3\]
rlabel metal2 97720 140952 97720 140952 0 A_all\[4\]
rlabel metal2 100856 140840 100856 140840 0 A_all\[5\]
rlabel metal2 93352 139846 93352 139846 0 A_all\[6\]
rlabel metal2 117544 143094 117544 143094 0 A_all\[7\]
rlabel metal2 118216 143878 118216 143878 0 A_all\[8\]
rlabel metal2 397110 259112 397110 259112 0 CEN_all
rlabel metal2 303464 551502 303464 551502 0 DAC_clk
rlabel metal2 313320 551558 313320 551558 0 DAC_d1
rlabel metal2 452872 499688 452872 499688 0 DAC_d2
rlabel metal2 308392 551446 308392 551446 0 DAC_le
rlabel metal2 145432 140742 145432 140742 0 D_all\[0\]
rlabel metal2 235032 139174 235032 139174 0 D_all\[1\]
rlabel metal2 233926 139048 233926 139048 0 D_all\[2\]
rlabel metal2 123368 143486 123368 143486 0 D_all\[3\]
rlabel metal2 122696 140112 122696 140112 0 D_all\[4\]
rlabel metal2 75544 140182 75544 140182 0 D_all\[5\]
rlabel metal2 74200 140518 74200 140518 0 D_all\[6\]
rlabel metal2 164584 142128 164584 142128 0 D_all\[7\]
rlabel metal2 106680 147350 106680 147350 0 GWEN_0
rlabel metal2 206584 142310 206584 142310 0 GWEN_1
rlabel metal2 138936 157906 138936 157906 0 GWEN_2
rlabel metal2 141624 157738 141624 157738 0 GWEN_3
rlabel metal2 144312 156058 144312 156058 0 GWEN_4
rlabel metal2 147000 159810 147000 159810 0 GWEN_5
rlabel metal3 307384 258776 307384 258776 0 GWEN_6
rlabel metal2 212184 212926 212184 212926 0 GWEN_7
rlabel metal2 143864 141750 143864 141750 0 Q0\[0\]
rlabel metal2 135688 141414 135688 141414 0 Q0\[1\]
rlabel metal2 133112 141582 133112 141582 0 Q0\[2\]
rlabel metal2 125048 142366 125048 142366 0 Q0\[3\]
rlabel metal2 149128 150472 149128 150472 0 Q0\[4\]
rlabel metal2 76104 143038 76104 143038 0 Q0\[5\]
rlabel metal2 73528 142254 73528 142254 0 Q0\[6\]
rlabel metal2 168504 155218 168504 155218 0 Q0\[7\]
rlabel metal2 171192 153538 171192 153538 0 Q1\[0\]
rlabel metal2 235704 141246 235704 141246 0 Q1\[1\]
rlabel metal2 233128 143094 233128 143094 0 Q1\[2\]
rlabel metal2 224952 141526 224952 141526 0 Q1\[3\]
rlabel metal2 184296 143486 184296 143486 0 Q1\[4\]
rlabel metal3 180376 152824 180376 152824 0 Q1\[5\]
rlabel metal2 187320 152866 187320 152866 0 Q1\[6\]
rlabel metal2 165368 141582 165368 141582 0 Q1\[7\]
rlabel metal2 192696 158578 192696 158578 0 Q2\[0\]
rlabel metal2 195384 158634 195384 158634 0 Q2\[1\]
rlabel metal2 333144 144830 333144 144830 0 Q2\[2\]
rlabel metal2 200760 157962 200760 157962 0 Q2\[3\]
rlabel metal2 284312 145670 284312 145670 0 Q2\[4\]
rlabel metal2 276136 141582 276136 141582 0 Q2\[5\]
rlabel metal2 208824 158746 208824 158746 0 Q2\[6\]
rlabel metal2 265384 143206 265384 143206 0 Q2\[7\]
rlabel metal2 214200 157794 214200 157794 0 Q3\[0\]
rlabel metal2 216888 158802 216888 158802 0 Q3\[1\]
rlabel metal2 219576 155218 219576 155218 0 Q3\[2\]
rlabel metal2 424984 145614 424984 145614 0 Q3\[3\]
rlabel metal2 384398 139048 384398 139048 0 Q3\[4\]
rlabel metal2 376152 142366 376152 142366 0 Q3\[5\]
rlabel metal2 373464 141526 373464 141526 0 Q3\[6\]
rlabel metal2 233016 152922 233016 152922 0 Q3\[7\]
rlabel metal2 543928 141358 543928 141358 0 Q4\[0\]
rlabel metal2 238392 152754 238392 152754 0 Q4\[1\]
rlabel metal2 241080 152810 241080 152810 0 Q4\[2\]
rlabel metal2 525000 141414 525000 141414 0 Q4\[3\]
rlabel metal2 261240 150528 261240 150528 0 Q4\[4\]
rlabel metal2 476056 143038 476056 143038 0 Q4\[5\]
rlabel metal2 258664 155960 258664 155960 0 Q4\[6\]
rlabel metal2 265496 153888 265496 153888 0 Q4\[7\]
rlabel metal2 257208 159754 257208 159754 0 Q5\[0\]
rlabel metal2 260456 158928 260456 158928 0 Q5\[1\]
rlabel metal2 262584 158970 262584 158970 0 Q5\[2\]
rlabel metal2 265272 158802 265272 158802 0 Q5\[3\]
rlabel metal2 308280 156632 308280 156632 0 Q5\[4\]
rlabel metal2 542920 158914 542920 158914 0 Q5\[5\]
rlabel metal2 545496 158858 545496 158858 0 Q5\[6\]
rlabel metal2 276024 158970 276024 158970 0 Q5\[7\]
rlabel metal2 216216 234822 216216 234822 0 Q6\[0\]
rlabel metal2 220248 211638 220248 211638 0 Q6\[1\]
rlabel metal2 432642 259112 432642 259112 0 Q6\[2\]
rlabel metal2 424578 259112 424578 259112 0 Q6\[3\]
rlabel metal2 232344 234430 232344 234430 0 Q6\[4\]
rlabel metal2 376152 260638 376152 260638 0 Q6\[5\]
rlabel metal2 373464 260806 373464 260806 0 Q6\[6\]
rlabel metal2 357112 240240 357112 240240 0 Q6\[7\]
rlabel metal2 248472 239974 248472 239974 0 Q7\[0\]
rlabel metal3 311640 275576 311640 275576 0 Q7\[1\]
rlabel metal2 256536 212982 256536 212982 0 Q7\[2\]
rlabel metal2 260568 216342 260568 216342 0 Q7\[3\]
rlabel metal2 264600 239078 264600 239078 0 Q7\[4\]
rlabel metal3 319984 266504 319984 266504 0 Q7\[5\]
rlabel metal2 350280 244664 350280 244664 0 Q7\[6\]
rlabel metal3 382872 275576 382872 275576 0 Q7\[7\]
rlabel metal4 289912 304971 289912 304971 0 RAM_end_addr\[0\]
rlabel metal4 475496 326415 475496 326415 0 RAM_end_addr\[10\]
rlabel metal4 476280 333883 476280 333883 0 RAM_end_addr\[11\]
rlabel metal3 435330 328552 435330 328552 0 RAM_end_addr\[12\]
rlabel metal4 475720 334869 475720 334869 0 RAM_end_addr\[13\]
rlabel metal4 475496 330637 475496 330637 0 RAM_end_addr\[14\]
rlabel metal4 475608 331805 475608 331805 0 RAM_end_addr\[15\]
rlabel metal4 475608 318153 475608 318153 0 RAM_end_addr\[1\]
rlabel metal4 473144 300048 473144 300048 0 RAM_end_addr\[2\]
rlabel metal4 472920 300440 472920 300440 0 RAM_end_addr\[3\]
rlabel metal4 283080 306535 283080 306535 0 RAM_end_addr\[4\]
rlabel metal4 53592 337819 53592 337819 0 RAM_end_addr\[5\]
rlabel metal2 476952 312760 476952 312760 0 RAM_end_addr\[6\]
rlabel metal4 54376 340873 54376 340873 0 RAM_end_addr\[7\]
rlabel metal4 53704 337225 53704 337225 0 RAM_end_addr\[8\]
rlabel metal2 476504 313208 476504 313208 0 RAM_end_addr\[9\]
rlabel metal4 78120 315630 78120 315630 0 RAM_start_addr\[0\]
rlabel metal4 54824 324589 54824 324589 0 RAM_start_addr\[10\]
rlabel metal4 475496 312945 475496 312945 0 RAM_start_addr\[11\]
rlabel metal4 55048 325753 55048 325753 0 RAM_start_addr\[12\]
rlabel metal4 475496 314651 475496 314651 0 RAM_start_addr\[13\]
rlabel metal4 475496 286303 475496 286303 0 RAM_start_addr\[14\]
rlabel metal2 476840 307104 476840 307104 0 RAM_start_addr\[15\]
rlabel metal4 476840 295685 476840 295685 0 RAM_start_addr\[1\]
rlabel metal4 54600 318133 54600 318133 0 RAM_start_addr\[2\]
rlabel metal4 54712 314944 54712 314944 0 RAM_start_addr\[3\]
rlabel metal4 69720 320220 69720 320220 0 RAM_start_addr\[4\]
rlabel metal4 54936 316456 54936 316456 0 RAM_start_addr\[5\]
rlabel metal4 475496 308185 475496 308185 0 RAM_start_addr\[6\]
rlabel metal4 53368 319963 53368 319963 0 RAM_start_addr\[7\]
rlabel metal4 53256 324775 53256 324775 0 RAM_start_addr\[8\]
rlabel metal4 53480 322207 53480 322207 0 RAM_start_addr\[9\]
rlabel metal2 284760 449736 284760 449736 0 RXD
rlabel metal2 194152 498274 194152 498274 0 TXD
rlabel metal2 144718 139048 144718 139048 0 WEN_all\[0\]
rlabel metal2 235032 142072 235032 142072 0 WEN_all\[1\]
rlabel metal2 235144 141792 235144 141792 0 WEN_all\[2\]
rlabel metal2 123690 139048 123690 139048 0 WEN_all\[3\]
rlabel metal2 186424 141624 186424 141624 0 WEN_all\[4\]
rlabel metal2 75096 140574 75096 140574 0 WEN_all\[5\]
rlabel metal2 74648 140630 74648 140630 0 WEN_all\[6\]
rlabel metal2 164472 140182 164472 140182 0 WEN_all\[7\]
rlabel metal2 71064 211414 71064 211414 0 WEb_ram
rlabel metal3 470680 452802 470680 452802 0 bus_addr\[0\]
rlabel metal3 214424 505778 214424 505778 0 bus_addr\[1\]
rlabel metal3 214998 508536 214998 508536 0 bus_addr\[2\]
rlabel metal4 468664 403869 468664 403869 0 bus_addr\[3\]
rlabel metal3 469210 477400 469210 477400 0 bus_addr\[4\]
rlabel metal2 169302 429912 169302 429912 0 bus_addr\[5\]
rlabel metal3 431536 549304 431536 549304 0 bus_cyc
rlabel metal4 474712 390768 474712 390768 0 bus_data_gpios\[0\]
rlabel metal4 472920 393232 472920 393232 0 bus_data_gpios\[1\]
rlabel metal4 454440 392392 454440 392392 0 bus_data_gpios\[2\]
rlabel metal4 474824 398104 474824 398104 0 bus_data_gpios\[3\]
rlabel metal4 452760 395304 452760 395304 0 bus_data_gpios\[4\]
rlabel metal3 363006 384776 363006 384776 0 bus_data_gpios\[5\]
rlabel metal4 449400 398216 449400 398216 0 bus_data_gpios\[6\]
rlabel metal4 451080 399672 451080 399672 0 bus_data_gpios\[7\]
rlabel metal3 470792 450296 470792 450296 0 bus_data_out\[0\]
rlabel metal3 469336 450408 469336 450408 0 bus_data_out\[1\]
rlabel metal3 470120 501242 470120 501242 0 bus_data_out\[2\]
rlabel metal3 214872 519638 214872 519638 0 bus_data_out\[3\]
rlabel metal3 214872 521794 214872 521794 0 bus_data_out\[4\]
rlabel metal3 216230 524664 216230 524664 0 bus_data_out\[5\]
rlabel metal3 469322 525784 469322 525784 0 bus_data_out\[6\]
rlabel metal3 471632 446824 471632 446824 0 bus_data_out\[7\]
rlabel metal2 171570 429912 171570 429912 0 bus_data_serial_ports\[0\]
rlabel metal3 216734 535416 216734 535416 0 bus_data_serial_ports\[1\]
rlabel metal3 215166 538104 215166 538104 0 bus_data_serial_ports\[2\]
rlabel metal3 215110 540792 215110 540792 0 bus_data_serial_ports\[3\]
rlabel metal3 215054 543480 215054 543480 0 bus_data_serial_ports\[4\]
rlabel metal3 216678 546168 216678 546168 0 bus_data_serial_ports\[5\]
rlabel metal3 215334 548856 215334 548856 0 bus_data_serial_ports\[6\]
rlabel metal2 190456 434630 190456 434630 0 bus_data_serial_ports\[7\]
rlabel metal4 387016 548968 387016 548968 0 bus_data_sid\[0\]
rlabel metal3 283206 392840 283206 392840 0 bus_data_sid\[1\]
rlabel metal3 348432 549304 348432 549304 0 bus_data_sid\[2\]
rlabel metal2 406952 550494 406952 550494 0 bus_data_sid\[3\]
rlabel metal3 281526 396872 281526 396872 0 bus_data_sid\[4\]
rlabel metal3 272286 398216 272286 398216 0 bus_data_sid\[5\]
rlabel metal2 421736 551670 421736 551670 0 bus_data_sid\[6\]
rlabel metal2 426664 551726 426664 551726 0 bus_data_sid\[7\]
rlabel metal4 249592 428456 249592 428456 0 bus_data_timers\[0\]
rlabel metal4 252280 428512 252280 428512 0 bus_data_timers\[1\]
rlabel metal2 254968 430430 254968 430430 0 bus_data_timers\[2\]
rlabel metal2 257656 430486 257656 430486 0 bus_data_timers\[3\]
rlabel metal4 260344 416175 260344 416175 0 bus_data_timers\[4\]
rlabel metal3 263368 429240 263368 429240 0 bus_data_timers\[5\]
rlabel metal3 266392 433384 266392 433384 0 bus_data_timers\[6\]
rlabel metal2 268590 429912 268590 429912 0 bus_data_timers\[7\]
rlabel metal2 517048 379498 517048 379498 0 bus_we_gpios
rlabel metal3 227248 452872 227248 452872 0 bus_we_serial_ports
rlabel metal2 289800 471520 289800 471520 0 bus_we_sid
rlabel metal2 244216 430374 244216 430374 0 bus_we_timers
rlabel metal4 60760 366511 60760 366511 0 cs_port\[0\]
rlabel via4 60760 367993 60760 367993 0 cs_port\[1\]
rlabel metal2 492632 343294 492632 343294 0 cs_port\[2\]
rlabel metal2 565320 142688 565320 142688 0 io_in[0]
rlabel metal3 593362 403592 593362 403592 0 io_in[10]
rlabel metal2 91000 431438 91000 431438 0 io_in[11]
rlabel metal2 93688 430094 93688 430094 0 io_in[12]
rlabel metal3 593082 522760 593082 522760 0 io_in[13]
rlabel metal2 99064 432110 99064 432110 0 io_in[14]
rlabel metal4 584696 590537 584696 590537 0 io_in[15]
rlabel metal2 518504 593306 518504 593306 0 io_in[16]
rlabel metal2 121800 502376 121800 502376 0 io_in[17]
rlabel metal2 386120 593026 386120 593026 0 io_in[18]
rlabel metal2 320152 593474 320152 593474 0 io_in[19]
rlabel metal3 593082 46984 593082 46984 0 io_in[1]
rlabel metal2 253960 592298 253960 592298 0 io_in[20]
rlabel metal2 187544 575498 187544 575498 0 io_in[21]
rlabel metal2 121352 583002 121352 583002 0 io_in[22]
rlabel metal2 55384 593138 55384 593138 0 io_in[23]
rlabel metal3 228270 587160 228270 587160 0 io_in[24]
rlabel metal3 2366 545048 2366 545048 0 io_in[25]
rlabel metal3 2310 502488 2310 502488 0 io_in[26]
rlabel metal3 2422 460152 2422 460152 0 io_in[27]
rlabel metal3 2534 418040 2534 418040 0 io_in[28]
rlabel metal3 2310 375704 2310 375704 0 io_in[29]
rlabel metal2 52024 296296 52024 296296 0 io_in[2]
rlabel metal3 2310 333144 2310 333144 0 io_in[30]
rlabel metal3 2702 290808 2702 290808 0 io_in[31]
rlabel via4 4200 248481 4200 248481 0 io_in[32]
rlabel metal3 2310 206360 2310 206360 0 io_in[33]
rlabel metal3 2310 164024 2310 164024 0 io_in[34]
rlabel metal2 21000 261576 21000 261576 0 io_in[37]
rlabel metal2 69496 430094 69496 430094 0 io_in[3]
rlabel metal3 593138 165928 593138 165928 0 io_in[4]
rlabel via4 74872 429371 74872 429371 0 io_in[5]
rlabel metal4 77560 431863 77560 431863 0 io_in[6]
rlabel metal4 590184 285041 590184 285041 0 io_in[7]
rlabel metal3 593082 324520 593082 324520 0 io_in[8]
rlabel metal2 279832 406224 279832 406224 0 io_in[9]
rlabel metal3 54936 300776 54936 300776 0 io_oeb[0]
rlabel metal3 593250 430136 593250 430136 0 io_oeb[10]
rlabel metal3 593250 469672 593250 469672 0 io_oeb[11]
rlabel metal4 478072 425275 478072 425275 0 io_oeb[12]
rlabel metal4 590184 548399 590184 548399 0 io_oeb[13]
rlabel metal4 52024 463512 52024 463512 0 io_oeb[14]
rlabel metal2 53704 460936 53704 460936 0 io_oeb[15]
rlabel metal2 55384 462448 55384 462448 0 io_oeb[16]
rlabel metal2 50344 465640 50344 465640 0 io_oeb[17]
rlabel metal3 200256 572152 200256 572152 0 io_oeb[18]
rlabel metal3 277032 590184 277032 590184 0 io_oeb[19]
rlabel metal3 593082 73416 593082 73416 0 io_oeb[1]
rlabel metal2 209832 593306 209832 593306 0 io_oeb[20]
rlabel metal2 143416 575442 143416 575442 0 io_oeb[21]
rlabel metal2 77336 580482 77336 580482 0 io_oeb[22]
rlabel metal2 490840 378826 490840 378826 0 io_oeb[23]
rlabel metal3 492856 380016 492856 380016 0 io_oeb[24]
rlabel metal3 2366 516600 2366 516600 0 io_oeb[25]
rlabel metal2 496888 379778 496888 379778 0 io_oeb[26]
rlabel metal4 498904 377747 498904 377747 0 io_oeb[27]
rlabel metal3 2422 389704 2422 389704 0 io_oeb[28]
rlabel metal3 2310 347480 2310 347480 0 io_oeb[29]
rlabel metal4 55272 233800 55272 233800 0 io_oeb[2]
rlabel metal3 2422 304920 2422 304920 0 io_oeb[30]
rlabel metal3 194670 262584 194670 262584 0 io_oeb[31]
rlabel metal3 2478 220472 2478 220472 0 io_oeb[32]
rlabel metal3 2366 178024 2366 178024 0 io_oeb[33]
rlabel metal3 2310 135800 2310 135800 0 io_oeb[34]
rlabel metal3 6510 93240 6510 93240 0 io_oeb[35]
rlabel metal2 185192 482314 185192 482314 0 io_oeb[36]
rlabel metal2 189672 483154 189672 483154 0 io_oeb[37]
rlabel metal3 59066 323624 59066 323624 0 io_oeb[3]
rlabel metal3 593138 192360 593138 192360 0 io_oeb[4]
rlabel metal3 593250 232008 593250 232008 0 io_oeb[5]
rlabel metal4 74760 299111 74760 299111 0 io_oeb[6]
rlabel metal3 593474 311080 593474 311080 0 io_oeb[7]
rlabel metal3 593362 350728 593362 350728 0 io_oeb[8]
rlabel metal4 53144 316189 53144 316189 0 io_oeb[9]
rlabel metal2 353640 145096 353640 145096 0 io_out[0]
rlabel metal4 76552 296550 76552 296550 0 io_out[10]
rlabel metal3 593138 456456 593138 456456 0 io_out[11]
rlabel metal3 593082 496104 593082 496104 0 io_out[12]
rlabel metal4 55384 431299 55384 431299 0 io_out[13]
rlabel metal4 50344 444136 50344 444136 0 io_out[14]
rlabel metal2 51912 446488 51912 446488 0 io_out[15]
rlabel metal2 496440 588938 496440 588938 0 io_out[16]
rlabel metal2 430248 580538 430248 580538 0 io_out[17]
rlabel metal3 210560 567000 210560 567000 0 io_out[18]
rlabel metal2 451304 520352 451304 520352 0 io_out[19]
rlabel metal4 567000 165648 567000 165648 0 io_out[1]
rlabel metal2 449400 512736 449400 512736 0 io_out[20]
rlabel metal2 165704 593250 165704 593250 0 io_out[21]
rlabel metal2 99512 593194 99512 593194 0 io_out[22]
rlabel metal2 451080 518336 451080 518336 0 io_out[23]
rlabel metal2 452760 503664 452760 503664 0 io_out[24]
rlabel metal3 2310 530824 2310 530824 0 io_out[25]
rlabel metal4 478408 415576 478408 415576 0 io_out[26]
rlabel metal3 2702 446040 2702 446040 0 io_out[27]
rlabel metal3 2366 403928 2366 403928 0 io_out[28]
rlabel metal3 2310 361592 2310 361592 0 io_out[29]
rlabel metal3 593250 99848 593250 99848 0 io_out[2]
rlabel metal3 2366 319032 2366 319032 0 io_out[30]
rlabel metal2 520002 429912 520002 429912 0 io_out[31]
rlabel metal3 2310 234584 2310 234584 0 io_out[32]
rlabel metal3 2422 192248 2422 192248 0 io_out[33]
rlabel metal2 524440 430038 524440 430038 0 io_out[34]
rlabel metal2 167272 473074 167272 473074 0 io_out[35]
rlabel metal3 3990 65240 3990 65240 0 io_out[36]
rlabel metal2 22680 245280 22680 245280 0 io_out[37]
rlabel metal2 568680 204456 568680 204456 0 io_out[3]
rlabel metal2 570360 227696 570360 227696 0 io_out[4]
rlabel metal3 593194 218792 593194 218792 0 io_out[5]
rlabel metal4 572040 263088 572040 263088 0 io_out[6]
rlabel metal4 55160 292807 55160 292807 0 io_out[7]
rlabel metal3 593418 337512 593418 337512 0 io_out[8]
rlabel metal4 590184 376815 590184 376815 0 io_out[9]
rlabel metal2 519064 379834 519064 379834 0 irq0
rlabel metal2 493528 448994 493528 448994 0 irq1
rlabel metal2 117880 431718 117880 431718 0 irq2
rlabel metal2 120568 449750 120568 449750 0 irq3
rlabel metal2 123256 431774 123256 431774 0 irq5
rlabel via4 521080 377927 521080 377927 0 irq6
rlabel metal3 490560 380128 490560 380128 0 irq7
rlabel metal2 215320 3150 215320 3150 0 la_data_out[0]
rlabel metal2 260344 76496 260344 76496 0 la_data_out[10]
rlabel metal2 277928 2310 277928 2310 0 la_data_out[11]
rlabel metal3 281680 5096 281680 5096 0 la_data_out[12]
rlabel metal3 288736 5096 288736 5096 0 la_data_out[13]
rlabel metal4 289800 161112 289800 161112 0 la_data_out[14]
rlabel metal3 297808 5096 297808 5096 0 la_data_out[15]
rlabel metal3 305704 4200 305704 4200 0 la_data_out[16]
rlabel metal2 312200 3206 312200 3206 0 la_data_out[17]
rlabel metal2 317912 3990 317912 3990 0 la_data_out[18]
rlabel metal3 323120 4200 323120 4200 0 la_data_out[19]
rlabel metal2 221032 3206 221032 3206 0 la_data_out[1]
rlabel metal2 329336 2310 329336 2310 0 la_data_out[20]
rlabel metal2 335272 2310 335272 2310 0 la_data_out[21]
rlabel metal3 271726 326984 271726 326984 0 la_data_out[22]
rlabel metal3 271614 328328 271614 328328 0 la_data_out[23]
rlabel metal2 352184 84630 352184 84630 0 la_data_out[24]
rlabel metal2 284760 250768 284760 250768 0 la_data_out[25]
rlabel metal2 350504 140784 350504 140784 0 la_data_out[26]
rlabel metal2 357000 130984 357000 130984 0 la_data_out[27]
rlabel metal2 375032 2646 375032 2646 0 la_data_out[28]
rlabel metal2 380744 2590 380744 2590 0 la_data_out[29]
rlabel metal2 226744 2254 226744 2254 0 la_data_out[2]
rlabel metal4 353640 164819 353640 164819 0 la_data_out[30]
rlabel metal3 284046 339080 284046 339080 0 la_data_out[31]
rlabel metal2 397880 2422 397880 2422 0 la_data_out[32]
rlabel metal2 403592 2478 403592 2478 0 la_data_out[33]
rlabel metal2 409304 3150 409304 3150 0 la_data_out[34]
rlabel metal2 415016 2366 415016 2366 0 la_data_out[35]
rlabel metal2 420728 8190 420728 8190 0 la_data_out[36]
rlabel metal4 284760 182392 284760 182392 0 la_data_out[37]
rlabel metal4 358680 173955 358680 173955 0 la_data_out[38]
rlabel metal4 355320 192795 355320 192795 0 la_data_out[39]
rlabel metal2 232456 2254 232456 2254 0 la_data_out[3]
rlabel metal2 443800 2310 443800 2310 0 la_data_out[40]
rlabel metal2 449288 76342 449288 76342 0 la_data_out[41]
rlabel metal2 455000 136038 455000 136038 0 la_data_out[42]
rlabel metal4 449512 196995 449512 196995 0 la_data_out[43]
rlabel metal4 452872 181151 452872 181151 0 la_data_out[44]
rlabel metal2 472136 2534 472136 2534 0 la_data_out[45]
rlabel metal2 477848 2478 477848 2478 0 la_data_out[46]
rlabel metal4 452760 181537 452760 181537 0 la_data_out[47]
rlabel metal3 271838 361928 271838 361928 0 la_data_out[48]
rlabel metal2 494984 2366 494984 2366 0 la_data_out[49]
rlabel metal2 238168 2534 238168 2534 0 la_data_out[4]
rlabel metal2 500696 3150 500696 3150 0 la_data_out[50]
rlabel metal4 451080 194565 451080 194565 0 la_data_out[51]
rlabel metal4 454552 202151 454552 202151 0 la_data_out[52]
rlabel metal2 517832 17430 517832 17430 0 la_data_out[53]
rlabel metal2 523544 2310 523544 2310 0 la_data_out[54]
rlabel metal4 451192 202095 451192 202095 0 la_data_out[55]
rlabel metal2 460152 227192 460152 227192 0 la_data_out[56]
rlabel metal2 540680 18270 540680 18270 0 la_data_out[57]
rlabel metal2 546616 2310 546616 2310 0 la_data_out[58]
rlabel metal2 468664 290136 468664 290136 0 la_data_out[59]
rlabel metal2 243880 2310 243880 2310 0 la_data_out[5]
rlabel metal2 477064 399168 477064 399168 0 la_data_out[60]
rlabel metal2 478632 399112 478632 399112 0 la_data_out[61]
rlabel metal2 478744 399056 478744 399056 0 la_data_out[62]
rlabel metal3 480088 427210 480088 427210 0 la_data_out[63]
rlabel metal3 264096 148680 264096 148680 0 la_data_out[6]
rlabel metal2 278936 229600 278936 229600 0 la_data_out[7]
rlabel metal2 260792 7350 260792 7350 0 la_data_out[8]
rlabel metal2 266728 2366 266728 2366 0 la_data_out[9]
rlabel metal4 475496 332343 475496 332343 0 last_addr\[0\]
rlabel metal4 475496 333331 475496 333331 0 last_addr\[1\]
rlabel metal2 476392 358904 476392 358904 0 last_addr\[2\]
rlabel metal2 209272 431270 209272 431270 0 last_addr\[3\]
rlabel metal2 212366 429912 212366 429912 0 last_addr\[4\]
rlabel metal2 214648 430206 214648 430206 0 last_addr\[5\]
rlabel metal4 475496 337551 475496 337551 0 last_addr\[6\]
rlabel metal2 220024 430318 220024 430318 0 last_addr\[7\]
rlabel metal2 512274 534968 512274 534968 0 pwm0
rlabel metal3 539742 399560 539742 399560 0 pwm1
rlabel metal2 546798 534968 546798 534968 0 pwm2
rlabel metal2 50008 350000 50008 350000 0 ram_bus_in\[0\]
rlabel metal2 48664 316120 48664 316120 0 ram_bus_in\[1\]
rlabel metal2 115416 249046 115416 249046 0 ram_bus_in\[2\]
rlabel metal2 119448 247422 119448 247422 0 ram_bus_in\[3\]
rlabel metal2 50232 324016 50232 324016 0 ram_bus_in\[4\]
rlabel metal3 60312 421666 60312 421666 0 ram_bus_in\[5\]
rlabel metal3 59234 423080 59234 423080 0 ram_bus_in\[6\]
rlabel metal3 60200 424130 60200 424130 0 ram_bus_in\[7\]
rlabel metal2 139608 246526 139608 246526 0 ram_enabled
rlabel metal2 143640 247366 143640 247366 0 requested_addr\[0\]
rlabel metal2 183960 212086 183960 212086 0 requested_addr\[10\]
rlabel metal2 187992 217126 187992 217126 0 requested_addr\[11\]
rlabel metal2 192024 246582 192024 246582 0 requested_addr\[12\]
rlabel metal2 196056 247478 196056 247478 0 requested_addr\[13\]
rlabel metal3 235424 283304 235424 283304 0 requested_addr\[14\]
rlabel metal3 237384 257880 237384 257880 0 requested_addr\[15\]
rlabel metal2 147672 246526 147672 246526 0 requested_addr\[1\]
rlabel metal3 211344 284872 211344 284872 0 requested_addr\[2\]
rlabel metal2 155736 213766 155736 213766 0 requested_addr\[3\]
rlabel metal2 159768 211246 159768 211246 0 requested_addr\[4\]
rlabel metal2 163800 216286 163800 216286 0 requested_addr\[5\]
rlabel metal2 167832 238182 167832 238182 0 requested_addr\[6\]
rlabel metal2 171864 211302 171864 211302 0 requested_addr\[7\]
rlabel metal2 175896 211358 175896 211358 0 requested_addr\[8\]
rlabel metal2 179928 211414 179928 211414 0 requested_addr\[9\]
rlabel metal4 212520 492184 212520 492184 0 reset
rlabel metal2 495992 343406 495992 343406 0 rom_bus_in\[0\]
rlabel metal2 499170 341880 499170 341880 0 rom_bus_in\[1\]
rlabel metal3 60312 407358 60312 407358 0 rom_bus_in\[2\]
rlabel metal3 189448 427560 189448 427560 0 rom_bus_in\[3\]
rlabel metal4 284984 386333 284984 386333 0 rom_bus_in\[4\]
rlabel metal3 176624 427224 176624 427224 0 rom_bus_in\[5\]
rlabel metal4 289800 386280 289800 386280 0 rom_bus_in\[6\]
rlabel metal4 281400 386460 281400 386460 0 rom_bus_in\[7\]
rlabel metal2 75096 211470 75096 211470 0 rom_bus_out\[0\]
rlabel metal2 53704 268464 53704 268464 0 rom_bus_out\[1\]
rlabel metal3 58184 354424 58184 354424 0 rom_bus_out\[2\]
rlabel metal2 48552 310128 48552 310128 0 rom_bus_out\[3\]
rlabel metal2 51800 341096 51800 341096 0 rom_bus_out\[4\]
rlabel metal2 95256 211246 95256 211246 0 rom_bus_out\[5\]
rlabel metal2 48440 329728 48440 329728 0 rom_bus_out\[6\]
rlabel metal2 50120 334656 50120 334656 0 rom_bus_out\[7\]
rlabel metal2 540568 448938 540568 448938 0 tmr0_clk
rlabel metal3 473984 537656 473984 537656 0 tmr0_o
rlabel metal2 549976 448882 549976 448882 0 tmr1_clk
rlabel metal2 495446 534968 495446 534968 0 tmr1_o
rlabel metal3 283206 372680 283206 372680 0 user_irq[0]
rlabel metal2 289800 320208 289800 320208 0 user_irq[1]
rlabel metal3 282422 375368 282422 375368 0 user_irq[2]
rlabel metal2 119336 140126 119336 140126 0 wb_clk_i
rlabel metal2 13384 2366 13384 2366 0 wb_rst_i
rlabel metal2 67256 287602 67256 287602 0 wbs_ack_o
rlabel metal2 23016 2254 23016 2254 0 wbs_adr_i[0]
rlabel metal4 148008 155344 148008 155344 0 wbs_adr_i[10]
rlabel metal2 93464 3990 93464 3990 0 wbs_adr_i[11]
rlabel metal2 99064 4046 99064 4046 0 wbs_adr_i[12]
rlabel metal3 153496 285656 153496 285656 0 wbs_adr_i[13]
rlabel metal2 159768 287896 159768 287896 0 wbs_adr_i[14]
rlabel metal2 116312 2254 116312 2254 0 wbs_adr_i[15]
rlabel metal2 122024 2534 122024 2534 0 wbs_adr_i[16]
rlabel metal2 148904 74200 148904 74200 0 wbs_adr_i[17]
rlabel metal4 143640 4424 143640 4424 0 wbs_adr_i[18]
rlabel metal2 139160 2758 139160 2758 0 wbs_adr_i[19]
rlabel metal2 30632 2646 30632 2646 0 wbs_adr_i[1]
rlabel metal2 144872 2590 144872 2590 0 wbs_adr_i[20]
rlabel metal3 173880 147224 173880 147224 0 wbs_adr_i[21]
rlabel metal2 208376 287882 208376 287882 0 wbs_adr_i[22]
rlabel metal2 162008 2422 162008 2422 0 wbs_adr_i[23]
rlabel metal2 167720 2310 167720 2310 0 wbs_adr_i[24]
rlabel metal2 173432 2142 173432 2142 0 wbs_adr_i[25]
rlabel metal2 231896 287896 231896 287896 0 wbs_adr_i[26]
rlabel metal3 238168 285656 238168 285656 0 wbs_adr_i[27]
rlabel metal2 190568 3990 190568 3990 0 wbs_adr_i[28]
rlabel metal2 196056 19110 196056 19110 0 wbs_adr_i[29]
rlabel metal2 38024 112350 38024 112350 0 wbs_adr_i[2]
rlabel metal3 256200 285656 256200 285656 0 wbs_adr_i[30]
rlabel metal3 260400 285880 260400 285880 0 wbs_adr_i[31]
rlabel metal2 45640 127470 45640 127470 0 wbs_adr_i[3]
rlabel metal2 53256 114870 53256 114870 0 wbs_adr_i[4]
rlabel metal3 82264 211176 82264 211176 0 wbs_adr_i[5]
rlabel metal3 62496 4200 62496 4200 0 wbs_adr_i[6]
rlabel metal2 70392 2310 70392 2310 0 wbs_adr_i[7]
rlabel metal2 123704 288274 123704 288274 0 wbs_adr_i[8]
rlabel metal2 82040 2310 82040 2310 0 wbs_adr_i[9]
rlabel metal2 24360 117600 24360 117600 0 wbs_cyc_i
rlabel metal2 24696 109046 24696 109046 0 wbs_dat_i[0]
rlabel metal2 137816 288162 137816 288162 0 wbs_dat_i[10]
rlabel metal2 143864 288330 143864 288330 0 wbs_dat_i[11]
rlabel metal2 101080 3150 101080 3150 0 wbs_dat_i[12]
rlabel metal3 155288 285656 155288 285656 0 wbs_dat_i[13]
rlabel metal2 162008 249746 162008 249746 0 wbs_dat_i[14]
rlabel metal2 118216 2310 118216 2310 0 wbs_dat_i[15]
rlabel metal2 123928 2366 123928 2366 0 wbs_dat_i[16]
rlabel metal2 129640 2198 129640 2198 0 wbs_dat_i[17]
rlabel metal3 185528 285656 185528 285656 0 wbs_dat_i[18]
rlabel metal2 141064 2646 141064 2646 0 wbs_dat_i[19]
rlabel metal2 32536 2366 32536 2366 0 wbs_dat_i[1]
rlabel metal2 146776 2702 146776 2702 0 wbs_dat_i[20]
rlabel metal2 152488 2366 152488 2366 0 wbs_dat_i[21]
rlabel metal2 210392 288498 210392 288498 0 wbs_dat_i[22]
rlabel metal2 163912 2478 163912 2478 0 wbs_dat_i[23]
rlabel metal2 169624 2366 169624 2366 0 wbs_dat_i[24]
rlabel metal2 175112 2534 175112 2534 0 wbs_dat_i[25]
rlabel metal2 234584 250474 234584 250474 0 wbs_dat_i[26]
rlabel metal2 186760 4046 186760 4046 0 wbs_dat_i[27]
rlabel metal2 192472 2366 192472 2366 0 wbs_dat_i[28]
rlabel metal2 252168 287896 252168 287896 0 wbs_dat_i[29]
rlabel metal2 44520 118776 44520 118776 0 wbs_dat_i[2]
rlabel metal3 258328 285656 258328 285656 0 wbs_dat_i[30]
rlabel metal3 262192 285768 262192 285768 0 wbs_dat_i[31]
rlabel metal2 47768 2310 47768 2310 0 wbs_dat_i[3]
rlabel metal2 55384 2702 55384 2702 0 wbs_dat_i[4]
rlabel metal3 60424 4312 60424 4312 0 wbs_dat_i[5]
rlabel metal3 63392 4424 63392 4424 0 wbs_dat_i[6]
rlabel metal2 119672 288330 119672 288330 0 wbs_dat_i[7]
rlabel metal2 78232 2310 78232 2310 0 wbs_dat_i[8]
rlabel metal4 121800 156296 121800 156296 0 wbs_dat_i[9]
rlabel metal2 26824 2310 26824 2310 0 wbs_dat_o[0]
rlabel metal3 139216 285656 139216 285656 0 wbs_dat_o[10]
rlabel metal2 145880 288050 145880 288050 0 wbs_dat_o[11]
rlabel metal2 102984 2310 102984 2310 0 wbs_dat_o[12]
rlabel metal2 108696 2310 108696 2310 0 wbs_dat_o[13]
rlabel metal2 114408 2310 114408 2310 0 wbs_dat_o[14]
rlabel metal2 170072 288498 170072 288498 0 wbs_dat_o[15]
rlabel metal2 125832 2422 125832 2422 0 wbs_dat_o[16]
rlabel metal2 131544 2254 131544 2254 0 wbs_dat_o[17]
rlabel metal2 188216 287882 188216 287882 0 wbs_dat_o[18]
rlabel metal2 194264 288386 194264 288386 0 wbs_dat_o[19]
rlabel metal2 51240 119448 51240 119448 0 wbs_dat_o[1]
rlabel metal2 148456 74550 148456 74550 0 wbs_dat_o[20]
rlabel metal4 167160 215488 167160 215488 0 wbs_dat_o[21]
rlabel metal2 212408 288330 212408 288330 0 wbs_dat_o[22]
rlabel metal2 165816 2254 165816 2254 0 wbs_dat_o[23]
rlabel metal3 171360 4200 171360 4200 0 wbs_dat_o[24]
rlabel metal3 229096 285768 229096 285768 0 wbs_dat_o[25]
rlabel metal2 236600 288274 236600 288274 0 wbs_dat_o[26]
rlabel metal2 188664 2254 188664 2254 0 wbs_dat_o[27]
rlabel metal2 194376 2310 194376 2310 0 wbs_dat_o[28]
rlabel metal4 258776 157920 258776 157920 0 wbs_dat_o[29]
rlabel metal2 91448 270634 91448 270634 0 wbs_dat_o[2]
rlabel metal3 260008 138936 260008 138936 0 wbs_dat_o[30]
rlabel metal2 211512 2478 211512 2478 0 wbs_dat_o[31]
rlabel metal3 97048 285656 97048 285656 0 wbs_dat_o[3]
rlabel metal3 59192 139384 59192 139384 0 wbs_dat_o[4]
rlabel metal3 61432 4088 61432 4088 0 wbs_dat_o[5]
rlabel metal2 68712 2366 68712 2366 0 wbs_dat_o[6]
rlabel metal2 74200 2254 74200 2254 0 wbs_dat_o[7]
rlabel metal4 123480 222600 123480 222600 0 wbs_dat_o[8]
rlabel metal2 85848 2366 85848 2366 0 wbs_dat_o[9]
rlabel metal2 71288 288442 71288 288442 0 wbs_stb_i
rlabel metal2 73304 288386 73304 288386 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
