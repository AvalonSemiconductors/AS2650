magic
tech gf180mcuC
magscale 1 5
timestamp 1695812890
<< obsm1 >>
rect 672 855 109312 78497
<< metal2 >>
rect 1176 79600 1232 80000
rect 2128 79600 2184 80000
rect 3080 79600 3136 80000
rect 4032 79600 4088 80000
rect 4984 79600 5040 80000
rect 5936 79600 5992 80000
rect 6888 79600 6944 80000
rect 7840 79600 7896 80000
rect 8792 79600 8848 80000
rect 9744 79600 9800 80000
rect 10696 79600 10752 80000
rect 11648 79600 11704 80000
rect 12600 79600 12656 80000
rect 13552 79600 13608 80000
rect 14504 79600 14560 80000
rect 15456 79600 15512 80000
rect 16408 79600 16464 80000
rect 17360 79600 17416 80000
rect 18312 79600 18368 80000
rect 19264 79600 19320 80000
rect 20216 79600 20272 80000
rect 21168 79600 21224 80000
rect 22120 79600 22176 80000
rect 23072 79600 23128 80000
rect 24024 79600 24080 80000
rect 24976 79600 25032 80000
rect 25928 79600 25984 80000
rect 26880 79600 26936 80000
rect 27832 79600 27888 80000
rect 28784 79600 28840 80000
rect 29736 79600 29792 80000
rect 30688 79600 30744 80000
rect 31640 79600 31696 80000
rect 32592 79600 32648 80000
rect 33544 79600 33600 80000
rect 34496 79600 34552 80000
rect 35448 79600 35504 80000
rect 36400 79600 36456 80000
rect 37352 79600 37408 80000
rect 38304 79600 38360 80000
rect 39256 79600 39312 80000
rect 40208 79600 40264 80000
rect 41160 79600 41216 80000
rect 42112 79600 42168 80000
rect 43064 79600 43120 80000
rect 44016 79600 44072 80000
rect 44968 79600 45024 80000
rect 45920 79600 45976 80000
rect 46872 79600 46928 80000
rect 47824 79600 47880 80000
rect 48776 79600 48832 80000
rect 49728 79600 49784 80000
rect 50680 79600 50736 80000
rect 51632 79600 51688 80000
rect 52584 79600 52640 80000
rect 53536 79600 53592 80000
rect 54488 79600 54544 80000
rect 55440 79600 55496 80000
rect 56392 79600 56448 80000
rect 57344 79600 57400 80000
rect 58296 79600 58352 80000
rect 59248 79600 59304 80000
rect 60200 79600 60256 80000
rect 61152 79600 61208 80000
rect 62104 79600 62160 80000
rect 63056 79600 63112 80000
rect 64008 79600 64064 80000
rect 64960 79600 65016 80000
rect 65912 79600 65968 80000
rect 66864 79600 66920 80000
rect 67816 79600 67872 80000
rect 68768 79600 68824 80000
rect 69720 79600 69776 80000
rect 70672 79600 70728 80000
rect 71624 79600 71680 80000
rect 72576 79600 72632 80000
rect 73528 79600 73584 80000
rect 74480 79600 74536 80000
rect 75432 79600 75488 80000
rect 76384 79600 76440 80000
rect 77336 79600 77392 80000
rect 78288 79600 78344 80000
rect 79240 79600 79296 80000
rect 80192 79600 80248 80000
rect 81144 79600 81200 80000
rect 82096 79600 82152 80000
rect 83048 79600 83104 80000
rect 84000 79600 84056 80000
rect 84952 79600 85008 80000
rect 85904 79600 85960 80000
rect 86856 79600 86912 80000
rect 87808 79600 87864 80000
rect 88760 79600 88816 80000
rect 89712 79600 89768 80000
rect 90664 79600 90720 80000
rect 91616 79600 91672 80000
rect 92568 79600 92624 80000
rect 93520 79600 93576 80000
rect 94472 79600 94528 80000
rect 95424 79600 95480 80000
rect 96376 79600 96432 80000
rect 97328 79600 97384 80000
rect 98280 79600 98336 80000
rect 99232 79600 99288 80000
rect 100184 79600 100240 80000
rect 101136 79600 101192 80000
rect 102088 79600 102144 80000
rect 103040 79600 103096 80000
rect 103992 79600 104048 80000
rect 104944 79600 105000 80000
rect 105896 79600 105952 80000
rect 106848 79600 106904 80000
rect 107800 79600 107856 80000
rect 108752 79600 108808 80000
rect 1176 0 1232 400
rect 2856 0 2912 400
rect 4536 0 4592 400
rect 6216 0 6272 400
rect 7896 0 7952 400
rect 9576 0 9632 400
rect 11256 0 11312 400
rect 12936 0 12992 400
rect 14616 0 14672 400
rect 16296 0 16352 400
rect 17976 0 18032 400
rect 19656 0 19712 400
rect 21336 0 21392 400
rect 23016 0 23072 400
rect 24696 0 24752 400
rect 26376 0 26432 400
rect 28056 0 28112 400
rect 29736 0 29792 400
rect 31416 0 31472 400
rect 33096 0 33152 400
rect 34776 0 34832 400
rect 36456 0 36512 400
rect 38136 0 38192 400
rect 39816 0 39872 400
rect 41496 0 41552 400
rect 43176 0 43232 400
rect 44856 0 44912 400
rect 46536 0 46592 400
rect 48216 0 48272 400
rect 49896 0 49952 400
rect 51576 0 51632 400
rect 53256 0 53312 400
rect 54936 0 54992 400
rect 56616 0 56672 400
rect 58296 0 58352 400
rect 59976 0 60032 400
rect 61656 0 61712 400
rect 63336 0 63392 400
rect 65016 0 65072 400
rect 66696 0 66752 400
rect 68376 0 68432 400
rect 70056 0 70112 400
rect 71736 0 71792 400
rect 73416 0 73472 400
rect 75096 0 75152 400
rect 76776 0 76832 400
rect 78456 0 78512 400
rect 80136 0 80192 400
rect 81816 0 81872 400
rect 83496 0 83552 400
rect 85176 0 85232 400
rect 86856 0 86912 400
rect 88536 0 88592 400
rect 90216 0 90272 400
rect 91896 0 91952 400
rect 93576 0 93632 400
rect 95256 0 95312 400
rect 96936 0 96992 400
rect 98616 0 98672 400
rect 100296 0 100352 400
rect 101976 0 102032 400
rect 103656 0 103712 400
rect 105336 0 105392 400
rect 107016 0 107072 400
rect 108696 0 108752 400
<< obsm2 >>
rect 742 79570 1146 79679
rect 1262 79570 2098 79679
rect 2214 79570 3050 79679
rect 3166 79570 4002 79679
rect 4118 79570 4954 79679
rect 5070 79570 5906 79679
rect 6022 79570 6858 79679
rect 6974 79570 7810 79679
rect 7926 79570 8762 79679
rect 8878 79570 9714 79679
rect 9830 79570 10666 79679
rect 10782 79570 11618 79679
rect 11734 79570 12570 79679
rect 12686 79570 13522 79679
rect 13638 79570 14474 79679
rect 14590 79570 15426 79679
rect 15542 79570 16378 79679
rect 16494 79570 17330 79679
rect 17446 79570 18282 79679
rect 18398 79570 19234 79679
rect 19350 79570 20186 79679
rect 20302 79570 21138 79679
rect 21254 79570 22090 79679
rect 22206 79570 23042 79679
rect 23158 79570 23994 79679
rect 24110 79570 24946 79679
rect 25062 79570 25898 79679
rect 26014 79570 26850 79679
rect 26966 79570 27802 79679
rect 27918 79570 28754 79679
rect 28870 79570 29706 79679
rect 29822 79570 30658 79679
rect 30774 79570 31610 79679
rect 31726 79570 32562 79679
rect 32678 79570 33514 79679
rect 33630 79570 34466 79679
rect 34582 79570 35418 79679
rect 35534 79570 36370 79679
rect 36486 79570 37322 79679
rect 37438 79570 38274 79679
rect 38390 79570 39226 79679
rect 39342 79570 40178 79679
rect 40294 79570 41130 79679
rect 41246 79570 42082 79679
rect 42198 79570 43034 79679
rect 43150 79570 43986 79679
rect 44102 79570 44938 79679
rect 45054 79570 45890 79679
rect 46006 79570 46842 79679
rect 46958 79570 47794 79679
rect 47910 79570 48746 79679
rect 48862 79570 49698 79679
rect 49814 79570 50650 79679
rect 50766 79570 51602 79679
rect 51718 79570 52554 79679
rect 52670 79570 53506 79679
rect 53622 79570 54458 79679
rect 54574 79570 55410 79679
rect 55526 79570 56362 79679
rect 56478 79570 57314 79679
rect 57430 79570 58266 79679
rect 58382 79570 59218 79679
rect 59334 79570 60170 79679
rect 60286 79570 61122 79679
rect 61238 79570 62074 79679
rect 62190 79570 63026 79679
rect 63142 79570 63978 79679
rect 64094 79570 64930 79679
rect 65046 79570 65882 79679
rect 65998 79570 66834 79679
rect 66950 79570 67786 79679
rect 67902 79570 68738 79679
rect 68854 79570 69690 79679
rect 69806 79570 70642 79679
rect 70758 79570 71594 79679
rect 71710 79570 72546 79679
rect 72662 79570 73498 79679
rect 73614 79570 74450 79679
rect 74566 79570 75402 79679
rect 75518 79570 76354 79679
rect 76470 79570 77306 79679
rect 77422 79570 78258 79679
rect 78374 79570 79210 79679
rect 79326 79570 80162 79679
rect 80278 79570 81114 79679
rect 81230 79570 82066 79679
rect 82182 79570 83018 79679
rect 83134 79570 83970 79679
rect 84086 79570 84922 79679
rect 85038 79570 85874 79679
rect 85990 79570 86826 79679
rect 86942 79570 87778 79679
rect 87894 79570 88730 79679
rect 88846 79570 89682 79679
rect 89798 79570 90634 79679
rect 90750 79570 91586 79679
rect 91702 79570 92538 79679
rect 92654 79570 93490 79679
rect 93606 79570 94442 79679
rect 94558 79570 95394 79679
rect 95510 79570 96346 79679
rect 96462 79570 97298 79679
rect 97414 79570 98250 79679
rect 98366 79570 99202 79679
rect 99318 79570 100154 79679
rect 100270 79570 101106 79679
rect 101222 79570 102058 79679
rect 102174 79570 103010 79679
rect 103126 79570 103962 79679
rect 104078 79570 104914 79679
rect 105030 79570 105866 79679
rect 105982 79570 106818 79679
rect 106934 79570 107770 79679
rect 107886 79570 108722 79679
rect 108838 79570 108906 79679
rect 742 430 108906 79570
rect 742 9 1146 430
rect 1262 9 2826 430
rect 2942 9 4506 430
rect 4622 9 6186 430
rect 6302 9 7866 430
rect 7982 9 9546 430
rect 9662 9 11226 430
rect 11342 9 12906 430
rect 13022 9 14586 430
rect 14702 9 16266 430
rect 16382 9 17946 430
rect 18062 9 19626 430
rect 19742 9 21306 430
rect 21422 9 22986 430
rect 23102 9 24666 430
rect 24782 9 26346 430
rect 26462 9 28026 430
rect 28142 9 29706 430
rect 29822 9 31386 430
rect 31502 9 33066 430
rect 33182 9 34746 430
rect 34862 9 36426 430
rect 36542 9 38106 430
rect 38222 9 39786 430
rect 39902 9 41466 430
rect 41582 9 43146 430
rect 43262 9 44826 430
rect 44942 9 46506 430
rect 46622 9 48186 430
rect 48302 9 49866 430
rect 49982 9 51546 430
rect 51662 9 53226 430
rect 53342 9 54906 430
rect 55022 9 56586 430
rect 56702 9 58266 430
rect 58382 9 59946 430
rect 60062 9 61626 430
rect 61742 9 63306 430
rect 63422 9 64986 430
rect 65102 9 66666 430
rect 66782 9 68346 430
rect 68462 9 70026 430
rect 70142 9 71706 430
rect 71822 9 73386 430
rect 73502 9 75066 430
rect 75182 9 76746 430
rect 76862 9 78426 430
rect 78542 9 80106 430
rect 80222 9 81786 430
rect 81902 9 83466 430
rect 83582 9 85146 430
rect 85262 9 86826 430
rect 86942 9 88506 430
rect 88622 9 90186 430
rect 90302 9 91866 430
rect 91982 9 93546 430
rect 93662 9 95226 430
rect 95342 9 96906 430
rect 97022 9 98586 430
rect 98702 9 100266 430
rect 100382 9 101946 430
rect 102062 9 103626 430
rect 103742 9 105306 430
rect 105422 9 106986 430
rect 107102 9 108666 430
rect 108782 9 108906 430
<< obsm3 >>
rect 737 14 102215 79674
<< metal4 >>
rect 2224 1538 2384 78430
rect 9904 1538 10064 78430
rect 17584 1538 17744 78430
rect 25264 1538 25424 78430
rect 32944 1538 33104 78430
rect 40624 1538 40784 78430
rect 48304 1538 48464 78430
rect 55984 1538 56144 78430
rect 63664 1538 63824 78430
rect 71344 1538 71504 78430
rect 79024 1538 79184 78430
rect 86704 1538 86864 78430
rect 94384 1538 94544 78430
rect 102064 1538 102224 78430
<< obsm4 >>
rect 4998 78460 80458 79343
rect 4998 1508 9874 78460
rect 10094 1508 17554 78460
rect 17774 1508 25234 78460
rect 25454 1508 32914 78460
rect 33134 1508 40594 78460
rect 40814 1508 48274 78460
rect 48494 1508 55954 78460
rect 56174 1508 63634 78460
rect 63854 1508 71314 78460
rect 71534 1508 78994 78460
rect 79214 1508 80458 78460
rect 4998 9 80458 1508
<< labels >>
rlabel metal2 s 1176 79600 1232 80000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 29736 79600 29792 80000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 32592 79600 32648 80000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 35448 79600 35504 80000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 38304 79600 38360 80000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 41160 79600 41216 80000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 44016 79600 44072 80000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 46872 79600 46928 80000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 49728 79600 49784 80000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 52584 79600 52640 80000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 55440 79600 55496 80000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4032 79600 4088 80000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 58296 79600 58352 80000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 61152 79600 61208 80000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 64008 79600 64064 80000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 66864 79600 66920 80000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 69720 79600 69776 80000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 72576 79600 72632 80000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 75432 79600 75488 80000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 78288 79600 78344 80000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 81144 79600 81200 80000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 84000 79600 84056 80000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6888 79600 6944 80000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 86856 79600 86912 80000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 89712 79600 89768 80000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 92568 79600 92624 80000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 95424 79600 95480 80000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 98280 79600 98336 80000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 101136 79600 101192 80000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 103992 79600 104048 80000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 106848 79600 106904 80000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9744 79600 9800 80000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 12600 79600 12656 80000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 15456 79600 15512 80000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 18312 79600 18368 80000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 21168 79600 21224 80000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 24024 79600 24080 80000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 26880 79600 26936 80000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2128 79600 2184 80000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 30688 79600 30744 80000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 33544 79600 33600 80000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 36400 79600 36456 80000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 39256 79600 39312 80000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 42112 79600 42168 80000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 44968 79600 45024 80000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 47824 79600 47880 80000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 50680 79600 50736 80000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 53536 79600 53592 80000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 56392 79600 56448 80000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 4984 79600 5040 80000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 59248 79600 59304 80000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 62104 79600 62160 80000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 64960 79600 65016 80000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 67816 79600 67872 80000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 70672 79600 70728 80000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 73528 79600 73584 80000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 76384 79600 76440 80000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 79240 79600 79296 80000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 82096 79600 82152 80000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 84952 79600 85008 80000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7840 79600 7896 80000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 87808 79600 87864 80000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 90664 79600 90720 80000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 93520 79600 93576 80000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 96376 79600 96432 80000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 99232 79600 99288 80000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 102088 79600 102144 80000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 104944 79600 105000 80000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 107800 79600 107856 80000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 10696 79600 10752 80000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 13552 79600 13608 80000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 16408 79600 16464 80000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 19264 79600 19320 80000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 22120 79600 22176 80000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 24976 79600 25032 80000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 27832 79600 27888 80000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3080 79600 3136 80000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 31640 79600 31696 80000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 34496 79600 34552 80000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 37352 79600 37408 80000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 40208 79600 40264 80000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 43064 79600 43120 80000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 45920 79600 45976 80000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 48776 79600 48832 80000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 51632 79600 51688 80000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 54488 79600 54544 80000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 57344 79600 57400 80000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5936 79600 5992 80000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 60200 79600 60256 80000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 63056 79600 63112 80000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 65912 79600 65968 80000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 68768 79600 68824 80000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 71624 79600 71680 80000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 74480 79600 74536 80000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 77336 79600 77392 80000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 80192 79600 80248 80000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 83048 79600 83104 80000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 85904 79600 85960 80000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8792 79600 8848 80000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 88760 79600 88816 80000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 91616 79600 91672 80000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 94472 79600 94528 80000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 97328 79600 97384 80000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 100184 79600 100240 80000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 103040 79600 103096 80000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 105896 79600 105952 80000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 108752 79600 108808 80000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 11648 79600 11704 80000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 14504 79600 14560 80000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 17360 79600 17416 80000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 20216 79600 20272 80000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 23072 79600 23128 80000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 25928 79600 25984 80000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 28784 79600 28840 80000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 2856 0 2912 400 6 la_data_out[0]
port 115 nsew signal output
rlabel metal2 s 19656 0 19712 400 6 la_data_out[10]
port 116 nsew signal output
rlabel metal2 s 21336 0 21392 400 6 la_data_out[11]
port 117 nsew signal output
rlabel metal2 s 23016 0 23072 400 6 la_data_out[12]
port 118 nsew signal output
rlabel metal2 s 24696 0 24752 400 6 la_data_out[13]
port 119 nsew signal output
rlabel metal2 s 26376 0 26432 400 6 la_data_out[14]
port 120 nsew signal output
rlabel metal2 s 28056 0 28112 400 6 la_data_out[15]
port 121 nsew signal output
rlabel metal2 s 29736 0 29792 400 6 la_data_out[16]
port 122 nsew signal output
rlabel metal2 s 31416 0 31472 400 6 la_data_out[17]
port 123 nsew signal output
rlabel metal2 s 33096 0 33152 400 6 la_data_out[18]
port 124 nsew signal output
rlabel metal2 s 34776 0 34832 400 6 la_data_out[19]
port 125 nsew signal output
rlabel metal2 s 4536 0 4592 400 6 la_data_out[1]
port 126 nsew signal output
rlabel metal2 s 36456 0 36512 400 6 la_data_out[20]
port 127 nsew signal output
rlabel metal2 s 38136 0 38192 400 6 la_data_out[21]
port 128 nsew signal output
rlabel metal2 s 39816 0 39872 400 6 la_data_out[22]
port 129 nsew signal output
rlabel metal2 s 41496 0 41552 400 6 la_data_out[23]
port 130 nsew signal output
rlabel metal2 s 43176 0 43232 400 6 la_data_out[24]
port 131 nsew signal output
rlabel metal2 s 44856 0 44912 400 6 la_data_out[25]
port 132 nsew signal output
rlabel metal2 s 46536 0 46592 400 6 la_data_out[26]
port 133 nsew signal output
rlabel metal2 s 48216 0 48272 400 6 la_data_out[27]
port 134 nsew signal output
rlabel metal2 s 49896 0 49952 400 6 la_data_out[28]
port 135 nsew signal output
rlabel metal2 s 51576 0 51632 400 6 la_data_out[29]
port 136 nsew signal output
rlabel metal2 s 6216 0 6272 400 6 la_data_out[2]
port 137 nsew signal output
rlabel metal2 s 53256 0 53312 400 6 la_data_out[30]
port 138 nsew signal output
rlabel metal2 s 54936 0 54992 400 6 la_data_out[31]
port 139 nsew signal output
rlabel metal2 s 56616 0 56672 400 6 la_data_out[32]
port 140 nsew signal output
rlabel metal2 s 58296 0 58352 400 6 la_data_out[33]
port 141 nsew signal output
rlabel metal2 s 59976 0 60032 400 6 la_data_out[34]
port 142 nsew signal output
rlabel metal2 s 61656 0 61712 400 6 la_data_out[35]
port 143 nsew signal output
rlabel metal2 s 63336 0 63392 400 6 la_data_out[36]
port 144 nsew signal output
rlabel metal2 s 65016 0 65072 400 6 la_data_out[37]
port 145 nsew signal output
rlabel metal2 s 66696 0 66752 400 6 la_data_out[38]
port 146 nsew signal output
rlabel metal2 s 68376 0 68432 400 6 la_data_out[39]
port 147 nsew signal output
rlabel metal2 s 7896 0 7952 400 6 la_data_out[3]
port 148 nsew signal output
rlabel metal2 s 70056 0 70112 400 6 la_data_out[40]
port 149 nsew signal output
rlabel metal2 s 71736 0 71792 400 6 la_data_out[41]
port 150 nsew signal output
rlabel metal2 s 73416 0 73472 400 6 la_data_out[42]
port 151 nsew signal output
rlabel metal2 s 75096 0 75152 400 6 la_data_out[43]
port 152 nsew signal output
rlabel metal2 s 76776 0 76832 400 6 la_data_out[44]
port 153 nsew signal output
rlabel metal2 s 78456 0 78512 400 6 la_data_out[45]
port 154 nsew signal output
rlabel metal2 s 80136 0 80192 400 6 la_data_out[46]
port 155 nsew signal output
rlabel metal2 s 81816 0 81872 400 6 la_data_out[47]
port 156 nsew signal output
rlabel metal2 s 83496 0 83552 400 6 la_data_out[48]
port 157 nsew signal output
rlabel metal2 s 85176 0 85232 400 6 la_data_out[49]
port 158 nsew signal output
rlabel metal2 s 9576 0 9632 400 6 la_data_out[4]
port 159 nsew signal output
rlabel metal2 s 86856 0 86912 400 6 la_data_out[50]
port 160 nsew signal output
rlabel metal2 s 88536 0 88592 400 6 la_data_out[51]
port 161 nsew signal output
rlabel metal2 s 90216 0 90272 400 6 la_data_out[52]
port 162 nsew signal output
rlabel metal2 s 91896 0 91952 400 6 la_data_out[53]
port 163 nsew signal output
rlabel metal2 s 93576 0 93632 400 6 la_data_out[54]
port 164 nsew signal output
rlabel metal2 s 95256 0 95312 400 6 la_data_out[55]
port 165 nsew signal output
rlabel metal2 s 96936 0 96992 400 6 la_data_out[56]
port 166 nsew signal output
rlabel metal2 s 98616 0 98672 400 6 la_data_out[57]
port 167 nsew signal output
rlabel metal2 s 100296 0 100352 400 6 la_data_out[58]
port 168 nsew signal output
rlabel metal2 s 101976 0 102032 400 6 la_data_out[59]
port 169 nsew signal output
rlabel metal2 s 11256 0 11312 400 6 la_data_out[5]
port 170 nsew signal output
rlabel metal2 s 103656 0 103712 400 6 la_data_out[60]
port 171 nsew signal output
rlabel metal2 s 105336 0 105392 400 6 la_data_out[61]
port 172 nsew signal output
rlabel metal2 s 107016 0 107072 400 6 la_data_out[62]
port 173 nsew signal output
rlabel metal2 s 108696 0 108752 400 6 la_data_out[63]
port 174 nsew signal output
rlabel metal2 s 12936 0 12992 400 6 la_data_out[6]
port 175 nsew signal output
rlabel metal2 s 14616 0 14672 400 6 la_data_out[7]
port 176 nsew signal output
rlabel metal2 s 16296 0 16352 400 6 la_data_out[8]
port 177 nsew signal output
rlabel metal2 s 17976 0 18032 400 6 la_data_out[9]
port 178 nsew signal output
rlabel metal4 s 2224 1538 2384 78430 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 78430 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 78430 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 78430 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 78430 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 78430 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 78430 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 78430 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 78430 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 78430 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 78430 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 78430 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 78430 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 78430 6 vss
port 180 nsew ground bidirectional
rlabel metal2 s 1176 0 1232 400 6 wb_clk_i
port 181 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17983344
string GDS_FILE /home/lucah/Desktop/AS2650/openlane/wrapped_as2650/runs/23_09_27_13_02/results/signoff/wrapped_as2650.magic.gds
string GDS_START 436660
<< end >>

