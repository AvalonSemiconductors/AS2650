magic
tech gf180mcuD
magscale 1 10
timestamp 1700712079
<< nwell >>
rect 1258 55257 298678 56096
rect 1258 55232 135821 55257
rect 1258 54503 131496 54528
rect 1258 53689 298678 54503
rect 1258 53664 191149 53689
rect 1258 52935 183309 52960
rect 1258 52096 298678 52935
rect 1258 50528 298678 51392
rect 1258 48960 298678 49824
rect 1258 47392 298678 48256
rect 1258 45824 298678 46688
rect 1258 44256 298678 45120
rect 1258 42688 298678 43552
rect 1258 41120 298678 41984
rect 1258 39552 298678 40416
rect 1258 37984 298678 38848
rect 1258 36416 298678 37280
rect 1258 34848 298678 35712
rect 1258 33280 298678 34144
rect 1258 31712 298678 32576
rect 1258 30144 298678 31008
rect 1258 28576 298678 29440
rect 1258 27008 298678 27872
rect 1258 25440 298678 26304
rect 1258 23872 298678 24736
rect 1258 22304 298678 23168
rect 1258 20736 298678 21600
rect 1258 19168 298678 20032
rect 1258 17600 298678 18464
rect 1258 16032 298678 16896
rect 1258 14464 298678 15328
rect 1258 12896 298678 13760
rect 1258 11328 298678 12192
rect 1258 9760 298678 10624
rect 1258 9031 192605 9056
rect 1258 8192 298678 9031
rect 1258 7463 185325 7488
rect 1258 6624 298678 7463
rect 1258 5895 183421 5920
rect 1258 5081 298678 5895
rect 1258 5056 182413 5081
rect 1258 4327 183421 4352
rect 1258 3513 298678 4327
rect 1258 3488 192381 3513
<< pwell >>
rect 1258 56096 298678 56534
rect 1258 54528 298678 55232
rect 1258 52960 298678 53664
rect 1258 51392 298678 52096
rect 1258 49824 298678 50528
rect 1258 48256 298678 48960
rect 1258 46688 298678 47392
rect 1258 45120 298678 45824
rect 1258 43552 298678 44256
rect 1258 41984 298678 42688
rect 1258 40416 298678 41120
rect 1258 38848 298678 39552
rect 1258 37280 298678 37984
rect 1258 35712 298678 36416
rect 1258 34144 298678 34848
rect 1258 32576 298678 33280
rect 1258 31008 298678 31712
rect 1258 29440 298678 30144
rect 1258 27872 298678 28576
rect 1258 26304 298678 27008
rect 1258 24736 298678 25440
rect 1258 23168 298678 23872
rect 1258 21600 298678 22304
rect 1258 20032 298678 20736
rect 1258 18464 298678 19168
rect 1258 16896 298678 17600
rect 1258 15328 298678 16032
rect 1258 13760 298678 14464
rect 1258 12192 298678 12896
rect 1258 10624 298678 11328
rect 1258 9056 298678 9760
rect 1258 7488 298678 8192
rect 1258 5920 298678 6624
rect 1258 4352 298678 5056
rect 1258 3050 298678 3488
<< obsm1 >>
rect 1344 3076 298592 57090
<< metal2 >>
rect 7392 59200 7504 60000
rect 12768 59200 12880 60000
rect 18144 59200 18256 60000
rect 23520 59200 23632 60000
rect 28896 59200 29008 60000
rect 34272 59200 34384 60000
rect 39648 59200 39760 60000
rect 45024 59200 45136 60000
rect 50400 59200 50512 60000
rect 55776 59200 55888 60000
rect 61152 59200 61264 60000
rect 66528 59200 66640 60000
rect 71904 59200 72016 60000
rect 77280 59200 77392 60000
rect 82656 59200 82768 60000
rect 88032 59200 88144 60000
rect 93408 59200 93520 60000
rect 98784 59200 98896 60000
rect 104160 59200 104272 60000
rect 109536 59200 109648 60000
rect 114912 59200 115024 60000
rect 120288 59200 120400 60000
rect 125664 59200 125776 60000
rect 131040 59200 131152 60000
rect 136416 59200 136528 60000
rect 141792 59200 141904 60000
rect 147168 59200 147280 60000
rect 152544 59200 152656 60000
rect 157920 59200 158032 60000
rect 163296 59200 163408 60000
rect 168672 59200 168784 60000
rect 174048 59200 174160 60000
rect 179424 59200 179536 60000
rect 184800 59200 184912 60000
rect 190176 59200 190288 60000
rect 195552 59200 195664 60000
rect 200928 59200 201040 60000
rect 206304 59200 206416 60000
rect 211680 59200 211792 60000
rect 217056 59200 217168 60000
rect 222432 59200 222544 60000
rect 227808 59200 227920 60000
rect 233184 59200 233296 60000
rect 238560 59200 238672 60000
rect 243936 59200 244048 60000
rect 249312 59200 249424 60000
rect 254688 59200 254800 60000
rect 260064 59200 260176 60000
rect 265440 59200 265552 60000
rect 270816 59200 270928 60000
rect 276192 59200 276304 60000
rect 281568 59200 281680 60000
rect 286944 59200 287056 60000
rect 292320 59200 292432 60000
rect 8288 0 8400 800
rect 11872 0 11984 800
rect 15456 0 15568 800
rect 19040 0 19152 800
rect 22624 0 22736 800
rect 26208 0 26320 800
rect 29792 0 29904 800
rect 33376 0 33488 800
rect 36960 0 37072 800
rect 40544 0 40656 800
rect 44128 0 44240 800
rect 47712 0 47824 800
rect 51296 0 51408 800
rect 54880 0 54992 800
rect 58464 0 58576 800
rect 62048 0 62160 800
rect 65632 0 65744 800
rect 69216 0 69328 800
rect 72800 0 72912 800
rect 76384 0 76496 800
rect 79968 0 80080 800
rect 83552 0 83664 800
rect 87136 0 87248 800
rect 90720 0 90832 800
rect 94304 0 94416 800
rect 97888 0 98000 800
rect 101472 0 101584 800
rect 105056 0 105168 800
rect 108640 0 108752 800
rect 112224 0 112336 800
rect 115808 0 115920 800
rect 119392 0 119504 800
rect 122976 0 123088 800
rect 126560 0 126672 800
rect 130144 0 130256 800
rect 133728 0 133840 800
rect 137312 0 137424 800
rect 140896 0 141008 800
rect 144480 0 144592 800
rect 148064 0 148176 800
rect 151648 0 151760 800
rect 155232 0 155344 800
rect 158816 0 158928 800
rect 162400 0 162512 800
rect 165984 0 166096 800
rect 169568 0 169680 800
rect 173152 0 173264 800
rect 176736 0 176848 800
rect 180320 0 180432 800
rect 183904 0 184016 800
rect 187488 0 187600 800
rect 191072 0 191184 800
rect 194656 0 194768 800
rect 198240 0 198352 800
rect 201824 0 201936 800
rect 205408 0 205520 800
rect 208992 0 209104 800
rect 212576 0 212688 800
rect 216160 0 216272 800
rect 219744 0 219856 800
rect 223328 0 223440 800
rect 226912 0 227024 800
rect 230496 0 230608 800
rect 234080 0 234192 800
rect 237664 0 237776 800
rect 241248 0 241360 800
rect 244832 0 244944 800
rect 248416 0 248528 800
rect 252000 0 252112 800
rect 255584 0 255696 800
rect 259168 0 259280 800
rect 262752 0 262864 800
rect 266336 0 266448 800
rect 269920 0 270032 800
rect 273504 0 273616 800
rect 277088 0 277200 800
rect 280672 0 280784 800
rect 284256 0 284368 800
rect 287840 0 287952 800
rect 291424 0 291536 800
<< obsm2 >>
rect 4476 59140 7332 59200
rect 7564 59140 12708 59200
rect 12940 59140 18084 59200
rect 18316 59140 23460 59200
rect 23692 59140 28836 59200
rect 29068 59140 34212 59200
rect 34444 59140 39588 59200
rect 39820 59140 44964 59200
rect 45196 59140 50340 59200
rect 50572 59140 55716 59200
rect 55948 59140 61092 59200
rect 61324 59140 66468 59200
rect 66700 59140 71844 59200
rect 72076 59140 77220 59200
rect 77452 59140 82596 59200
rect 82828 59140 87972 59200
rect 88204 59140 93348 59200
rect 93580 59140 98724 59200
rect 98956 59140 104100 59200
rect 104332 59140 109476 59200
rect 109708 59140 114852 59200
rect 115084 59140 120228 59200
rect 120460 59140 125604 59200
rect 125836 59140 130980 59200
rect 131212 59140 136356 59200
rect 136588 59140 141732 59200
rect 141964 59140 147108 59200
rect 147340 59140 152484 59200
rect 152716 59140 157860 59200
rect 158092 59140 163236 59200
rect 163468 59140 168612 59200
rect 168844 59140 173988 59200
rect 174220 59140 179364 59200
rect 179596 59140 184740 59200
rect 184972 59140 190116 59200
rect 190348 59140 195492 59200
rect 195724 59140 200868 59200
rect 201100 59140 206244 59200
rect 206476 59140 211620 59200
rect 211852 59140 216996 59200
rect 217228 59140 222372 59200
rect 222604 59140 227748 59200
rect 227980 59140 233124 59200
rect 233356 59140 238500 59200
rect 238732 59140 243876 59200
rect 244108 59140 249252 59200
rect 249484 59140 254628 59200
rect 254860 59140 260004 59200
rect 260236 59140 265380 59200
rect 265612 59140 270756 59200
rect 270988 59140 276132 59200
rect 276364 59140 281508 59200
rect 281740 59140 286884 59200
rect 287116 59140 292260 59200
rect 292492 59140 296580 59200
rect 4476 860 296580 59140
rect 4476 700 8228 860
rect 8460 700 11812 860
rect 12044 700 15396 860
rect 15628 700 18980 860
rect 19212 700 22564 860
rect 22796 700 26148 860
rect 26380 700 29732 860
rect 29964 700 33316 860
rect 33548 700 36900 860
rect 37132 700 40484 860
rect 40716 700 44068 860
rect 44300 700 47652 860
rect 47884 700 51236 860
rect 51468 700 54820 860
rect 55052 700 58404 860
rect 58636 700 61988 860
rect 62220 700 65572 860
rect 65804 700 69156 860
rect 69388 700 72740 860
rect 72972 700 76324 860
rect 76556 700 79908 860
rect 80140 700 83492 860
rect 83724 700 87076 860
rect 87308 700 90660 860
rect 90892 700 94244 860
rect 94476 700 97828 860
rect 98060 700 101412 860
rect 101644 700 104996 860
rect 105228 700 108580 860
rect 108812 700 112164 860
rect 112396 700 115748 860
rect 115980 700 119332 860
rect 119564 700 122916 860
rect 123148 700 126500 860
rect 126732 700 130084 860
rect 130316 700 133668 860
rect 133900 700 137252 860
rect 137484 700 140836 860
rect 141068 700 144420 860
rect 144652 700 148004 860
rect 148236 700 151588 860
rect 151820 700 155172 860
rect 155404 700 158756 860
rect 158988 700 162340 860
rect 162572 700 165924 860
rect 166156 700 169508 860
rect 169740 700 173092 860
rect 173324 700 176676 860
rect 176908 700 180260 860
rect 180492 700 183844 860
rect 184076 700 187428 860
rect 187660 700 191012 860
rect 191244 700 194596 860
rect 194828 700 198180 860
rect 198412 700 201764 860
rect 201996 700 205348 860
rect 205580 700 208932 860
rect 209164 700 212516 860
rect 212748 700 216100 860
rect 216332 700 219684 860
rect 219916 700 223268 860
rect 223500 700 226852 860
rect 227084 700 230436 860
rect 230668 700 234020 860
rect 234252 700 237604 860
rect 237836 700 241188 860
rect 241420 700 244772 860
rect 245004 700 248356 860
rect 248588 700 251940 860
rect 252172 700 255524 860
rect 255756 700 259108 860
rect 259340 700 262692 860
rect 262924 700 266276 860
rect 266508 700 269860 860
rect 270092 700 273444 860
rect 273676 700 277028 860
rect 277260 700 280612 860
rect 280844 700 284196 860
rect 284428 700 287780 860
rect 288012 700 291364 860
rect 291596 700 296580 860
<< obsm3 >>
rect 4466 1036 296590 56476
<< metal4 >>
rect 4448 3076 4768 56508
rect 19808 3076 20128 56508
rect 35168 3076 35488 56508
rect 50528 3076 50848 56508
rect 65888 3076 66208 56508
rect 81248 3076 81568 56508
rect 96608 3076 96928 56508
rect 111968 3076 112288 56508
rect 127328 3076 127648 56508
rect 142688 3076 143008 56508
rect 158048 3076 158368 56508
rect 173408 3076 173728 56508
rect 188768 3076 189088 56508
rect 204128 3076 204448 56508
rect 219488 3076 219808 56508
rect 234848 3076 235168 56508
rect 250208 3076 250528 56508
rect 265568 3076 265888 56508
rect 280928 3076 281248 56508
rect 296288 3076 296608 56508
<< obsm4 >>
rect 217084 4498 219428 10510
rect 219868 4498 220836 10510
<< labels >>
rlabel metal2 s 40544 0 40656 800 6 A_all[0]
port 1 nsew signal output
rlabel metal2 s 44128 0 44240 800 6 A_all[1]
port 2 nsew signal output
rlabel metal2 s 47712 0 47824 800 6 A_all[2]
port 3 nsew signal output
rlabel metal2 s 51296 0 51408 800 6 A_all[3]
port 4 nsew signal output
rlabel metal2 s 54880 0 54992 800 6 A_all[4]
port 5 nsew signal output
rlabel metal2 s 58464 0 58576 800 6 A_all[5]
port 6 nsew signal output
rlabel metal2 s 62048 0 62160 800 6 A_all[6]
port 7 nsew signal output
rlabel metal2 s 65632 0 65744 800 6 A_all[7]
port 8 nsew signal output
rlabel metal2 s 69216 0 69328 800 6 A_all[8]
port 9 nsew signal output
rlabel metal2 s 8288 0 8400 800 6 CEN_all
port 10 nsew signal output
rlabel metal2 s 72800 0 72912 800 6 D_all[0]
port 11 nsew signal output
rlabel metal2 s 76384 0 76496 800 6 D_all[1]
port 12 nsew signal output
rlabel metal2 s 79968 0 80080 800 6 D_all[2]
port 13 nsew signal output
rlabel metal2 s 83552 0 83664 800 6 D_all[3]
port 14 nsew signal output
rlabel metal2 s 87136 0 87248 800 6 D_all[4]
port 15 nsew signal output
rlabel metal2 s 90720 0 90832 800 6 D_all[5]
port 16 nsew signal output
rlabel metal2 s 94304 0 94416 800 6 D_all[6]
port 17 nsew signal output
rlabel metal2 s 97888 0 98000 800 6 D_all[7]
port 18 nsew signal output
rlabel metal2 s 101472 0 101584 800 6 GWEN_0
port 19 nsew signal output
rlabel metal2 s 105056 0 105168 800 6 GWEN_1
port 20 nsew signal output
rlabel metal2 s 108640 0 108752 800 6 GWEN_2
port 21 nsew signal output
rlabel metal2 s 112224 0 112336 800 6 GWEN_3
port 22 nsew signal output
rlabel metal2 s 115808 0 115920 800 6 GWEN_4
port 23 nsew signal output
rlabel metal2 s 119392 0 119504 800 6 GWEN_5
port 24 nsew signal output
rlabel metal2 s 200928 59200 201040 60000 6 GWEN_6
port 25 nsew signal output
rlabel metal2 s 206304 59200 206416 60000 6 GWEN_7
port 26 nsew signal output
rlabel metal2 s 122976 0 123088 800 6 Q0[0]
port 27 nsew signal input
rlabel metal2 s 126560 0 126672 800 6 Q0[1]
port 28 nsew signal input
rlabel metal2 s 130144 0 130256 800 6 Q0[2]
port 29 nsew signal input
rlabel metal2 s 133728 0 133840 800 6 Q0[3]
port 30 nsew signal input
rlabel metal2 s 137312 0 137424 800 6 Q0[4]
port 31 nsew signal input
rlabel metal2 s 140896 0 141008 800 6 Q0[5]
port 32 nsew signal input
rlabel metal2 s 144480 0 144592 800 6 Q0[6]
port 33 nsew signal input
rlabel metal2 s 148064 0 148176 800 6 Q0[7]
port 34 nsew signal input
rlabel metal2 s 151648 0 151760 800 6 Q1[0]
port 35 nsew signal input
rlabel metal2 s 155232 0 155344 800 6 Q1[1]
port 36 nsew signal input
rlabel metal2 s 158816 0 158928 800 6 Q1[2]
port 37 nsew signal input
rlabel metal2 s 162400 0 162512 800 6 Q1[3]
port 38 nsew signal input
rlabel metal2 s 165984 0 166096 800 6 Q1[4]
port 39 nsew signal input
rlabel metal2 s 169568 0 169680 800 6 Q1[5]
port 40 nsew signal input
rlabel metal2 s 173152 0 173264 800 6 Q1[6]
port 41 nsew signal input
rlabel metal2 s 176736 0 176848 800 6 Q1[7]
port 42 nsew signal input
rlabel metal2 s 180320 0 180432 800 6 Q2[0]
port 43 nsew signal input
rlabel metal2 s 183904 0 184016 800 6 Q2[1]
port 44 nsew signal input
rlabel metal2 s 187488 0 187600 800 6 Q2[2]
port 45 nsew signal input
rlabel metal2 s 191072 0 191184 800 6 Q2[3]
port 46 nsew signal input
rlabel metal2 s 194656 0 194768 800 6 Q2[4]
port 47 nsew signal input
rlabel metal2 s 198240 0 198352 800 6 Q2[5]
port 48 nsew signal input
rlabel metal2 s 201824 0 201936 800 6 Q2[6]
port 49 nsew signal input
rlabel metal2 s 205408 0 205520 800 6 Q2[7]
port 50 nsew signal input
rlabel metal2 s 208992 0 209104 800 6 Q3[0]
port 51 nsew signal input
rlabel metal2 s 212576 0 212688 800 6 Q3[1]
port 52 nsew signal input
rlabel metal2 s 216160 0 216272 800 6 Q3[2]
port 53 nsew signal input
rlabel metal2 s 219744 0 219856 800 6 Q3[3]
port 54 nsew signal input
rlabel metal2 s 223328 0 223440 800 6 Q3[4]
port 55 nsew signal input
rlabel metal2 s 226912 0 227024 800 6 Q3[5]
port 56 nsew signal input
rlabel metal2 s 230496 0 230608 800 6 Q3[6]
port 57 nsew signal input
rlabel metal2 s 234080 0 234192 800 6 Q3[7]
port 58 nsew signal input
rlabel metal2 s 237664 0 237776 800 6 Q4[0]
port 59 nsew signal input
rlabel metal2 s 241248 0 241360 800 6 Q4[1]
port 60 nsew signal input
rlabel metal2 s 244832 0 244944 800 6 Q4[2]
port 61 nsew signal input
rlabel metal2 s 248416 0 248528 800 6 Q4[3]
port 62 nsew signal input
rlabel metal2 s 252000 0 252112 800 6 Q4[4]
port 63 nsew signal input
rlabel metal2 s 255584 0 255696 800 6 Q4[5]
port 64 nsew signal input
rlabel metal2 s 259168 0 259280 800 6 Q4[6]
port 65 nsew signal input
rlabel metal2 s 262752 0 262864 800 6 Q4[7]
port 66 nsew signal input
rlabel metal2 s 266336 0 266448 800 6 Q5[0]
port 67 nsew signal input
rlabel metal2 s 269920 0 270032 800 6 Q5[1]
port 68 nsew signal input
rlabel metal2 s 273504 0 273616 800 6 Q5[2]
port 69 nsew signal input
rlabel metal2 s 277088 0 277200 800 6 Q5[3]
port 70 nsew signal input
rlabel metal2 s 280672 0 280784 800 6 Q5[4]
port 71 nsew signal input
rlabel metal2 s 284256 0 284368 800 6 Q5[5]
port 72 nsew signal input
rlabel metal2 s 287840 0 287952 800 6 Q5[6]
port 73 nsew signal input
rlabel metal2 s 291424 0 291536 800 6 Q5[7]
port 74 nsew signal input
rlabel metal2 s 211680 59200 211792 60000 6 Q6[0]
port 75 nsew signal input
rlabel metal2 s 217056 59200 217168 60000 6 Q6[1]
port 76 nsew signal input
rlabel metal2 s 222432 59200 222544 60000 6 Q6[2]
port 77 nsew signal input
rlabel metal2 s 227808 59200 227920 60000 6 Q6[3]
port 78 nsew signal input
rlabel metal2 s 233184 59200 233296 60000 6 Q6[4]
port 79 nsew signal input
rlabel metal2 s 238560 59200 238672 60000 6 Q6[5]
port 80 nsew signal input
rlabel metal2 s 243936 59200 244048 60000 6 Q6[6]
port 81 nsew signal input
rlabel metal2 s 249312 59200 249424 60000 6 Q6[7]
port 82 nsew signal input
rlabel metal2 s 254688 59200 254800 60000 6 Q7[0]
port 83 nsew signal input
rlabel metal2 s 260064 59200 260176 60000 6 Q7[1]
port 84 nsew signal input
rlabel metal2 s 265440 59200 265552 60000 6 Q7[2]
port 85 nsew signal input
rlabel metal2 s 270816 59200 270928 60000 6 Q7[3]
port 86 nsew signal input
rlabel metal2 s 276192 59200 276304 60000 6 Q7[4]
port 87 nsew signal input
rlabel metal2 s 281568 59200 281680 60000 6 Q7[5]
port 88 nsew signal input
rlabel metal2 s 286944 59200 287056 60000 6 Q7[6]
port 89 nsew signal input
rlabel metal2 s 292320 59200 292432 60000 6 Q7[7]
port 90 nsew signal input
rlabel metal2 s 11872 0 11984 800 6 WEN_all[0]
port 91 nsew signal output
rlabel metal2 s 15456 0 15568 800 6 WEN_all[1]
port 92 nsew signal output
rlabel metal2 s 19040 0 19152 800 6 WEN_all[2]
port 93 nsew signal output
rlabel metal2 s 22624 0 22736 800 6 WEN_all[3]
port 94 nsew signal output
rlabel metal2 s 26208 0 26320 800 6 WEN_all[4]
port 95 nsew signal output
rlabel metal2 s 29792 0 29904 800 6 WEN_all[5]
port 96 nsew signal output
rlabel metal2 s 33376 0 33488 800 6 WEN_all[6]
port 97 nsew signal output
rlabel metal2 s 36960 0 37072 800 6 WEN_all[7]
port 98 nsew signal output
rlabel metal2 s 18144 59200 18256 60000 6 WEb_raw
port 99 nsew signal input
rlabel metal2 s 23520 59200 23632 60000 6 bus_in[0]
port 100 nsew signal input
rlabel metal2 s 28896 59200 29008 60000 6 bus_in[1]
port 101 nsew signal input
rlabel metal2 s 34272 59200 34384 60000 6 bus_in[2]
port 102 nsew signal input
rlabel metal2 s 39648 59200 39760 60000 6 bus_in[3]
port 103 nsew signal input
rlabel metal2 s 45024 59200 45136 60000 6 bus_in[4]
port 104 nsew signal input
rlabel metal2 s 50400 59200 50512 60000 6 bus_in[5]
port 105 nsew signal input
rlabel metal2 s 55776 59200 55888 60000 6 bus_in[6]
port 106 nsew signal input
rlabel metal2 s 61152 59200 61264 60000 6 bus_in[7]
port 107 nsew signal input
rlabel metal2 s 66528 59200 66640 60000 6 bus_out[0]
port 108 nsew signal output
rlabel metal2 s 71904 59200 72016 60000 6 bus_out[1]
port 109 nsew signal output
rlabel metal2 s 77280 59200 77392 60000 6 bus_out[2]
port 110 nsew signal output
rlabel metal2 s 82656 59200 82768 60000 6 bus_out[3]
port 111 nsew signal output
rlabel metal2 s 88032 59200 88144 60000 6 bus_out[4]
port 112 nsew signal output
rlabel metal2 s 93408 59200 93520 60000 6 bus_out[5]
port 113 nsew signal output
rlabel metal2 s 98784 59200 98896 60000 6 bus_out[6]
port 114 nsew signal output
rlabel metal2 s 104160 59200 104272 60000 6 bus_out[7]
port 115 nsew signal output
rlabel metal2 s 109536 59200 109648 60000 6 ram_enabled
port 116 nsew signal input
rlabel metal2 s 114912 59200 115024 60000 6 requested_addr[0]
port 117 nsew signal input
rlabel metal2 s 168672 59200 168784 60000 6 requested_addr[10]
port 118 nsew signal input
rlabel metal2 s 174048 59200 174160 60000 6 requested_addr[11]
port 119 nsew signal input
rlabel metal2 s 179424 59200 179536 60000 6 requested_addr[12]
port 120 nsew signal input
rlabel metal2 s 184800 59200 184912 60000 6 requested_addr[13]
port 121 nsew signal input
rlabel metal2 s 190176 59200 190288 60000 6 requested_addr[14]
port 122 nsew signal input
rlabel metal2 s 195552 59200 195664 60000 6 requested_addr[15]
port 123 nsew signal input
rlabel metal2 s 120288 59200 120400 60000 6 requested_addr[1]
port 124 nsew signal input
rlabel metal2 s 125664 59200 125776 60000 6 requested_addr[2]
port 125 nsew signal input
rlabel metal2 s 131040 59200 131152 60000 6 requested_addr[3]
port 126 nsew signal input
rlabel metal2 s 136416 59200 136528 60000 6 requested_addr[4]
port 127 nsew signal input
rlabel metal2 s 141792 59200 141904 60000 6 requested_addr[5]
port 128 nsew signal input
rlabel metal2 s 147168 59200 147280 60000 6 requested_addr[6]
port 129 nsew signal input
rlabel metal2 s 152544 59200 152656 60000 6 requested_addr[7]
port 130 nsew signal input
rlabel metal2 s 157920 59200 158032 60000 6 requested_addr[8]
port 131 nsew signal input
rlabel metal2 s 163296 59200 163408 60000 6 requested_addr[9]
port 132 nsew signal input
rlabel metal2 s 12768 59200 12880 60000 6 rst
port 133 nsew signal input
rlabel metal4 s 4448 3076 4768 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 250208 3076 250528 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 280928 3076 281248 56508 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 234848 3076 235168 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 265568 3076 265888 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 296288 3076 296608 56508 6 vss
port 135 nsew ground bidirectional
rlabel metal2 s 7392 59200 7504 60000 6 wb_clk_i
port 136 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 300000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1912456
string GDS_FILE /run/media/tholin/d9eb5833-69bc-462f-98fb-b7c5c019399b/AS2650/openlane/ram_controller/runs/23_11_23_04_59/results/signoff/ram_controller.magic.gds
string GDS_START 184362
<< end >>

