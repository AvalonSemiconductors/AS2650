// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[13] ;
 wire \as2650.pc[14] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire net89;
 wire clknet_leaf_0_wb_clk_i;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net90;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net91;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net92;
 wire net93;
 wire net78;
 wire net83;
 wire net79;
 wire net80;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net81;
 wire net82;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_1_1_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;
 wire clknet_opt_2_1_wb_clk_i;
 wire clknet_opt_3_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4300_ (.I(net26),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4301_ (.I(\as2650.ins_reg[0] ),
    .Z(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4302_ (.I(_3882_),
    .Z(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4303_ (.I(_3883_),
    .ZN(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4304_ (.I(_3884_),
    .Z(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4305_ (.I(\as2650.psl[4] ),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4306_ (.I(_3886_),
    .Z(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4307_ (.I(_3887_),
    .Z(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4308_ (.I(_3888_),
    .Z(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4309_ (.I(_3889_),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4310_ (.I(\as2650.ins_reg[0] ),
    .Z(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4311_ (.I(\as2650.ins_reg[1] ),
    .Z(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4312_ (.A1(_3891_),
    .A2(_3892_),
    .ZN(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4313_ (.I(_3893_),
    .Z(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4314_ (.I(_3894_),
    .Z(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4315_ (.I(_3895_),
    .Z(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4316_ (.A1(_3890_),
    .A2(_3896_),
    .ZN(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4317_ (.I(_3897_),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4318_ (.I(\as2650.ins_reg[4] ),
    .Z(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4319_ (.I(_3899_),
    .Z(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4320_ (.I(_3900_),
    .Z(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4321_ (.I(\as2650.halted ),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4322_ (.I(net10),
    .ZN(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4323_ (.A1(_3902_),
    .A2(_3903_),
    .ZN(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4324_ (.I(_3904_),
    .Z(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4325_ (.A1(_3901_),
    .A2(_3905_),
    .ZN(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4326_ (.I(\as2650.cycle[7] ),
    .Z(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4327_ (.A1(\as2650.cycle[3] ),
    .A2(\as2650.cycle[2] ),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4328_ (.I(_3908_),
    .Z(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4329_ (.A1(\as2650.cycle[5] ),
    .A2(\as2650.cycle[4] ),
    .ZN(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4330_ (.A1(\as2650.cycle[6] ),
    .A2(_3910_),
    .Z(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4331_ (.I(\as2650.cycle[1] ),
    .Z(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4332_ (.I(\as2650.cycle[0] ),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4333_ (.A1(_3912_),
    .A2(_3913_),
    .ZN(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4334_ (.A1(_3909_),
    .A2(_3911_),
    .A3(_3914_),
    .Z(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4335_ (.I(_3915_),
    .Z(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4336_ (.A1(_3907_),
    .A2(_3916_),
    .ZN(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4337_ (.I(\as2650.addr_buff[6] ),
    .Z(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4338_ (.I(\as2650.addr_buff[5] ),
    .Z(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4339_ (.A1(_3918_),
    .A2(_3919_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4340_ (.A1(\as2650.addr_buff[7] ),
    .A2(_3920_),
    .Z(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4341_ (.A1(_3917_),
    .A2(_3921_),
    .ZN(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4342_ (.A1(_3906_),
    .A2(_3922_),
    .Z(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4343_ (.A1(_3898_),
    .A2(_3923_),
    .ZN(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4344_ (.I(_3890_),
    .Z(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4345_ (.A1(_3925_),
    .A2(_3904_),
    .ZN(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4346_ (.I(_3908_),
    .Z(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4347_ (.A1(\as2650.cycle[5] ),
    .A2(\as2650.cycle[4] ),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4348_ (.A1(\as2650.cycle[7] ),
    .A2(\as2650.cycle[6] ),
    .A3(_3928_),
    .ZN(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4349_ (.I(\as2650.cycle[1] ),
    .ZN(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4350_ (.A1(_3930_),
    .A2(\as2650.cycle[0] ),
    .ZN(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4351_ (.A1(_3929_),
    .A2(_3931_),
    .Z(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4352_ (.A1(_3927_),
    .A2(_3932_),
    .Z(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4353_ (.I(_3933_),
    .Z(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4354_ (.A1(_3926_),
    .A2(_3934_),
    .ZN(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4355_ (.I(_3896_),
    .Z(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4356_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .ZN(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4357_ (.I(_3937_),
    .Z(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4358_ (.I(_3938_),
    .Z(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4359_ (.I(_3939_),
    .Z(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4360_ (.I(_3940_),
    .Z(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4361_ (.I(_3899_),
    .ZN(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4362_ (.I(_3942_),
    .Z(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4363_ (.I(\as2650.ins_reg[5] ),
    .Z(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4364_ (.I(\as2650.ins_reg[6] ),
    .Z(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4365_ (.I(_3945_),
    .ZN(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4366_ (.I(\as2650.ins_reg[7] ),
    .Z(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4367_ (.I(_3947_),
    .ZN(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4368_ (.I(_3948_),
    .Z(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4369_ (.A1(_3944_),
    .A2(_3946_),
    .A3(_3949_),
    .ZN(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4370_ (.A1(_3943_),
    .A2(_3950_),
    .Z(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4371_ (.A1(_3941_),
    .A2(_3951_),
    .ZN(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4372_ (.A1(_3935_),
    .A2(_3936_),
    .A3(_3952_),
    .ZN(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4373_ (.I(_3953_),
    .Z(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4374_ (.I(\as2650.cycle[0] ),
    .Z(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4375_ (.A1(_3912_),
    .A2(_3955_),
    .A3(_3927_),
    .A4(_3929_),
    .ZN(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4376_ (.I(\as2650.ins_reg[2] ),
    .Z(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4377_ (.I(_3899_),
    .Z(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4378_ (.A1(_3958_),
    .A2(_3944_),
    .ZN(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4379_ (.A1(_3957_),
    .A2(_3959_),
    .ZN(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4380_ (.A1(_3949_),
    .A2(_3960_),
    .ZN(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4381_ (.A1(_3956_),
    .A2(_3961_),
    .ZN(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4382_ (.I(\as2650.ins_reg[3] ),
    .Z(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4383_ (.A1(_3963_),
    .A2(_3904_),
    .ZN(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4384_ (.I(_3964_),
    .Z(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4385_ (.A1(_3897_),
    .A2(_3962_),
    .A3(_3965_),
    .ZN(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4386_ (.I(_3966_),
    .Z(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4387_ (.I(_3967_),
    .ZN(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4388_ (.I(_3925_),
    .Z(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4389_ (.A1(_3969_),
    .A2(_3936_),
    .Z(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4390_ (.I(_3907_),
    .Z(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4391_ (.I(_3909_),
    .Z(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4392_ (.I(_3914_),
    .Z(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4393_ (.A1(_3972_),
    .A2(_3911_),
    .A3(_3973_),
    .ZN(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4394_ (.A1(_3971_),
    .A2(_3974_),
    .Z(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4395_ (.I(\as2650.idx_ctrl[1] ),
    .ZN(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4396_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4397_ (.A1(_3976_),
    .A2(_3977_),
    .ZN(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4398_ (.A1(_3906_),
    .A2(_3978_),
    .ZN(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4399_ (.A1(_3970_),
    .A2(_3975_),
    .A3(_3979_),
    .ZN(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4400_ (.A1(_3954_),
    .A2(_3968_),
    .A3(_3980_),
    .ZN(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4401_ (.I(_3929_),
    .Z(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4402_ (.A1(_3912_),
    .A2(\as2650.cycle[0] ),
    .ZN(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4403_ (.I(\as2650.cycle[2] ),
    .ZN(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4404_ (.A1(\as2650.cycle[3] ),
    .A2(_3984_),
    .ZN(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4405_ (.A1(_3983_),
    .A2(_3985_),
    .Z(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4406_ (.A1(_3982_),
    .A2(_3986_),
    .ZN(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4407_ (.A1(_3901_),
    .A2(_3987_),
    .ZN(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4408_ (.A1(\as2650.ins_reg[5] ),
    .A2(_3945_),
    .A3(_3947_),
    .ZN(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4409_ (.I(_3989_),
    .Z(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4410_ (.I(_3940_),
    .Z(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4411_ (.A1(_3936_),
    .A2(_3991_),
    .A3(_3978_),
    .ZN(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4412_ (.A1(_3988_),
    .A2(_3990_),
    .A3(_3992_),
    .ZN(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4413_ (.I(_3993_),
    .Z(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4414_ (.I(_3901_),
    .Z(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4415_ (.I(_3945_),
    .Z(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4416_ (.I(_3996_),
    .Z(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4417_ (.I(_3997_),
    .Z(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4418_ (.I(_3883_),
    .Z(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4419_ (.I(_3892_),
    .Z(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4420_ (.A1(_3999_),
    .A2(_4000_),
    .Z(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4421_ (.I(_4001_),
    .Z(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4422_ (.I(_4002_),
    .Z(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4423_ (.I(\as2650.ins_reg[3] ),
    .ZN(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4424_ (.I(_4004_),
    .Z(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4425_ (.I(_4005_),
    .Z(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4426_ (.A1(_3927_),
    .A2(_3932_),
    .ZN(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4427_ (.I(_4007_),
    .Z(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4428_ (.I(_4008_),
    .Z(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4429_ (.A1(_4006_),
    .A2(_4009_),
    .ZN(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4430_ (.A1(_3995_),
    .A2(_3998_),
    .A3(_4003_),
    .A4(_4010_),
    .ZN(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4431_ (.A1(_3994_),
    .A2(_4011_),
    .ZN(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4432_ (.A1(_3926_),
    .A2(_4012_),
    .ZN(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4433_ (.I(_3933_),
    .Z(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4434_ (.I(_4014_),
    .Z(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4435_ (.I(\as2650.ins_reg[5] ),
    .ZN(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4436_ (.A1(\as2650.ins_reg[4] ),
    .A2(\as2650.ins_reg[6] ),
    .A3(\as2650.ins_reg[7] ),
    .Z(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4437_ (.A1(_4016_),
    .A2(_4017_),
    .ZN(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4438_ (.A1(_3957_),
    .A2(_4018_),
    .ZN(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4439_ (.I(_4019_),
    .Z(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4440_ (.A1(_4015_),
    .A2(_3898_),
    .A3(_3965_),
    .A4(_4020_),
    .Z(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4441_ (.I(_4021_),
    .Z(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4442_ (.A1(_3926_),
    .A2(_4014_),
    .Z(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4443_ (.I(_4002_),
    .Z(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4444_ (.I(\as2650.ins_reg[2] ),
    .ZN(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4445_ (.I(\as2650.ins_reg[5] ),
    .Z(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4446_ (.A1(_3996_),
    .A2(_3949_),
    .ZN(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4447_ (.A1(_4026_),
    .A2(_4027_),
    .ZN(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4448_ (.A1(_4025_),
    .A2(_3900_),
    .A3(_4028_),
    .ZN(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4449_ (.A1(_3963_),
    .A2(_4029_),
    .ZN(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4450_ (.A1(_4023_),
    .A2(_4024_),
    .A3(_4030_),
    .Z(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4451_ (.I(_4031_),
    .Z(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4452_ (.A1(_4022_),
    .A2(_4032_),
    .ZN(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4453_ (.A1(_3924_),
    .A2(_3981_),
    .A3(_4013_),
    .A4(_4033_),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4454_ (.A1(_3885_),
    .A2(_4034_),
    .ZN(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4455_ (.I(_3969_),
    .Z(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4456_ (.I(_3905_),
    .Z(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4457_ (.A1(_4036_),
    .A2(_4037_),
    .A3(_3994_),
    .ZN(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4458_ (.I(_4038_),
    .Z(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4459_ (.A1(_3906_),
    .A2(_3922_),
    .ZN(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4460_ (.A1(_3970_),
    .A2(_4040_),
    .ZN(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4461_ (.I(_4041_),
    .Z(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4462_ (.I(_4042_),
    .Z(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4463_ (.A1(_3891_),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4464_ (.I(_3887_),
    .Z(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4465_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_4045_),
    .Z(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4466_ (.A1(_4044_),
    .A2(_4046_),
    .ZN(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4467_ (.I(\as2650.r0[0] ),
    .Z(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4468_ (.I(_4048_),
    .Z(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4469_ (.I(_4049_),
    .Z(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4470_ (.A1(\as2650.ins_reg[0] ),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4471_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123[0][0] ),
    .I2(\as2650.r123_2[1][0] ),
    .I3(\as2650.r123_2[0][0] ),
    .S0(_3891_),
    .S1(_4045_),
    .Z(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4472_ (.A1(_4050_),
    .A2(_3893_),
    .B1(_4051_),
    .B2(_4052_),
    .ZN(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4473_ (.A1(_4047_),
    .A2(_4053_),
    .Z(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4474_ (.I(_4054_),
    .Z(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4475_ (.I(\as2650.addr_buff[5] ),
    .ZN(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4476_ (.A1(_3918_),
    .A2(_4056_),
    .ZN(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4477_ (.I(\as2650.addr_buff[6] ),
    .ZN(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4478_ (.A1(_4058_),
    .A2(_3919_),
    .ZN(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4479_ (.A1(_4057_),
    .A2(_4059_),
    .ZN(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4480_ (.A1(_4055_),
    .A2(_4060_),
    .Z(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4481_ (.I(_4061_),
    .Z(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4482_ (.I(_4050_),
    .Z(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4483_ (.I(_4063_),
    .ZN(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4484_ (.I(_3953_),
    .Z(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4485_ (.I(_4065_),
    .Z(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4486_ (.I(_3954_),
    .Z(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4487_ (.I(net5),
    .Z(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4488_ (.I(_4068_),
    .Z(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4489_ (.I(_4069_),
    .Z(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4490_ (.I(_3966_),
    .Z(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4491_ (.I(_4071_),
    .Z(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4492_ (.A1(_4023_),
    .A2(_4024_),
    .A3(_4030_),
    .ZN(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4493_ (.I(_4073_),
    .Z(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4494_ (.I(_4054_),
    .Z(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4495_ (.A1(_4017_),
    .A2(_4075_),
    .Z(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4496_ (.A1(_3967_),
    .A2(_4076_),
    .ZN(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4497_ (.A1(_4070_),
    .A2(_4072_),
    .B(_4074_),
    .C(_4077_),
    .ZN(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4498_ (.I(_4031_),
    .Z(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4499_ (.I(_4044_),
    .Z(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4500_ (.I(_4045_),
    .Z(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4501_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_4081_),
    .Z(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4502_ (.A1(_4080_),
    .A2(_4082_),
    .ZN(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4503_ (.I(_4083_),
    .Z(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4504_ (.I(\as2650.r0[1] ),
    .Z(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4505_ (.I(_4085_),
    .Z(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4506_ (.I(_4051_),
    .Z(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4507_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123[0][1] ),
    .I2(\as2650.r123_2[1][1] ),
    .I3(\as2650.r123_2[0][1] ),
    .S0(_3882_),
    .S1(_4081_),
    .Z(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4508_ (.A1(_4086_),
    .A2(_3894_),
    .B1(_4087_),
    .B2(_4088_),
    .ZN(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4509_ (.I(_4089_),
    .Z(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4510_ (.A1(_4084_),
    .A2(_4090_),
    .ZN(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4511_ (.I(_4091_),
    .Z(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4512_ (.I(_4021_),
    .Z(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4513_ (.A1(_4079_),
    .A2(_4092_),
    .B(_4093_),
    .ZN(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4514_ (.I(\as2650.psl[3] ),
    .Z(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4515_ (.I(\as2650.r0[7] ),
    .Z(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4516_ (.I(_4096_),
    .Z(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4517_ (.A1(_4097_),
    .A2(_3896_),
    .ZN(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4518_ (.I(_4080_),
    .Z(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4519_ (.I(_4099_),
    .Z(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4520_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_3889_),
    .Z(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4521_ (.A1(_4100_),
    .A2(_4101_),
    .ZN(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4522_ (.I(_4087_),
    .Z(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4523_ (.I0(\as2650.r123[1][7] ),
    .I1(\as2650.r123[0][7] ),
    .I2(\as2650.r123_2[1][7] ),
    .I3(\as2650.r123_2[0][7] ),
    .S0(_3999_),
    .S1(_3890_),
    .Z(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4524_ (.A1(_4103_),
    .A2(_4104_),
    .ZN(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4525_ (.A1(_4098_),
    .A2(_4102_),
    .A3(_4105_),
    .ZN(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4526_ (.I(_4106_),
    .Z(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4527_ (.I(\as2650.carry ),
    .ZN(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4528_ (.A1(\as2650.psl[3] ),
    .A2(_4108_),
    .ZN(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4529_ (.A1(_4095_),
    .A2(_4107_),
    .B(_4109_),
    .ZN(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4530_ (.I(_4021_),
    .Z(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4531_ (.A1(_4078_),
    .A2(_4094_),
    .B1(_4110_),
    .B2(_4111_),
    .ZN(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4532_ (.A1(_4067_),
    .A2(_4112_),
    .ZN(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4533_ (.I(_4041_),
    .Z(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4534_ (.A1(_4064_),
    .A2(_4066_),
    .B(_4113_),
    .C(_4114_),
    .ZN(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4535_ (.I(_3980_),
    .Z(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4536_ (.A1(_4043_),
    .A2(_4062_),
    .B(_4115_),
    .C(_4116_),
    .ZN(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4537_ (.I(_3974_),
    .Z(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4538_ (.A1(_3971_),
    .A2(_4118_),
    .ZN(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4539_ (.I(_3958_),
    .Z(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4540_ (.I(_4120_),
    .Z(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4541_ (.I(_4121_),
    .Z(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4542_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4543_ (.A1(_4122_),
    .A2(_3905_),
    .A3(_4123_),
    .ZN(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4544_ (.A1(_3898_),
    .A2(_4119_),
    .A3(_4124_),
    .ZN(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4545_ (.I(_4125_),
    .Z(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4546_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_3977_),
    .ZN(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4547_ (.A1(_3976_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4548_ (.A1(_4127_),
    .A2(_4128_),
    .ZN(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4549_ (.A1(_4055_),
    .A2(_4129_),
    .Z(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4550_ (.I(_4130_),
    .Z(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4551_ (.A1(_4126_),
    .A2(_4131_),
    .ZN(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4552_ (.A1(_4117_),
    .A2(_4132_),
    .ZN(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4553_ (.I(_4047_),
    .Z(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4554_ (.I(_4053_),
    .Z(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4555_ (.I(\as2650.holding_reg[0] ),
    .ZN(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4556_ (.A1(_4134_),
    .A2(_4135_),
    .B(_4136_),
    .ZN(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4557_ (.I(_4136_),
    .Z(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4558_ (.I(_4134_),
    .Z(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4559_ (.I(_4135_),
    .Z(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4560_ (.A1(_4138_),
    .A2(_4139_),
    .A3(_4140_),
    .Z(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4561_ (.A1(_4137_),
    .A2(_4141_),
    .ZN(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4562_ (.I(_4026_),
    .Z(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4563_ (.I(_3947_),
    .Z(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4564_ (.A1(_3997_),
    .A2(_4144_),
    .ZN(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4565_ (.A1(_4143_),
    .A2(_4145_),
    .Z(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4566_ (.I(_4146_),
    .Z(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4567_ (.I(_4028_),
    .Z(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4568_ (.A1(_4103_),
    .A2(_4052_),
    .Z(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4569_ (.A1(_4100_),
    .A2(_4046_),
    .Z(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4570_ (.A1(_4064_),
    .A2(_4001_),
    .ZN(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4571_ (.A1(_4149_),
    .A2(_4150_),
    .A3(_4151_),
    .B(\as2650.holding_reg[0] ),
    .ZN(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4572_ (.A1(_4148_),
    .A2(_4152_),
    .B(_4146_),
    .ZN(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4573_ (.I(_4143_),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4574_ (.A1(_3996_),
    .A2(_3948_),
    .ZN(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4575_ (.I(_4155_),
    .Z(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4576_ (.A1(_4154_),
    .A2(_4156_),
    .ZN(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4577_ (.A1(_4109_),
    .A2(_4142_),
    .Z(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4578_ (.A1(_3946_),
    .A2(_4144_),
    .ZN(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4579_ (.A1(_4026_),
    .A2(_4159_),
    .ZN(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4580_ (.A1(\as2650.psl[3] ),
    .A2(\as2650.carry ),
    .ZN(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4581_ (.I(_4161_),
    .ZN(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4582_ (.A1(_4162_),
    .A2(_4142_),
    .Z(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4583_ (.I(_4016_),
    .Z(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(_4025_),
    .A2(_4004_),
    .ZN(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4585_ (.I(_4165_),
    .Z(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4586_ (.A1(_4138_),
    .A2(_4166_),
    .ZN(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4587_ (.A1(_4139_),
    .A2(_4140_),
    .B(_3938_),
    .ZN(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4588_ (.A1(_4167_),
    .A2(_4168_),
    .Z(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4589_ (.I(_4144_),
    .Z(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4590_ (.A1(_3946_),
    .A2(_4170_),
    .ZN(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4591_ (.I(_4171_),
    .Z(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4592_ (.A1(_4164_),
    .A2(_4169_),
    .B(_4172_),
    .ZN(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4593_ (.I(_3941_),
    .Z(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4594_ (.I(_4159_),
    .Z(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4595_ (.I(_4175_),
    .Z(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4596_ (.A1(_3941_),
    .A2(_4075_),
    .ZN(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4597_ (.A1(\as2650.holding_reg[0] ),
    .A2(_4174_),
    .B(_4176_),
    .C(_4177_),
    .ZN(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4598_ (.A1(_4173_),
    .A2(_4178_),
    .ZN(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4599_ (.A1(_4160_),
    .A2(_4163_),
    .B(_4179_),
    .ZN(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4600_ (.A1(_4157_),
    .A2(_4158_),
    .B(_4180_),
    .ZN(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4601_ (.A1(_4142_),
    .A2(_4147_),
    .B1(_4153_),
    .B2(_4181_),
    .ZN(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4602_ (.I(_4182_),
    .Z(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4603_ (.A1(_4039_),
    .A2(_4183_),
    .ZN(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4604_ (.A1(_4039_),
    .A2(_4133_),
    .B(_4184_),
    .ZN(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4605_ (.I(net10),
    .Z(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4606_ (.I(_4186_),
    .Z(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4607_ (.I(_4165_),
    .Z(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4608_ (.I(_4188_),
    .Z(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4609_ (.I(_4189_),
    .Z(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4610_ (.A1(_4002_),
    .A2(_4190_),
    .ZN(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4611_ (.I(_4026_),
    .Z(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4612_ (.A1(_3958_),
    .A2(_4155_),
    .ZN(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4613_ (.I(_4193_),
    .Z(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4614_ (.A1(_4192_),
    .A2(_4194_),
    .ZN(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4615_ (.A1(_4191_),
    .A2(_4195_),
    .ZN(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4616_ (.I(_4196_),
    .Z(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4617_ (.A1(_3935_),
    .A2(_4197_),
    .ZN(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4618_ (.I(_4198_),
    .Z(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4619_ (.I(_3999_),
    .Z(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4620_ (.I(_4200_),
    .Z(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4621_ (.I(_4201_),
    .Z(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4622_ (.A1(_4170_),
    .A2(_3959_),
    .ZN(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4623_ (.I(_3957_),
    .Z(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4624_ (.A1(_4204_),
    .A2(_3956_),
    .ZN(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4625_ (.A1(_4203_),
    .A2(_3964_),
    .A3(_4205_),
    .ZN(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4626_ (.A1(_3970_),
    .A2(_4206_),
    .ZN(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4627_ (.A1(_3953_),
    .A2(_4021_),
    .A3(_4031_),
    .A4(_4207_),
    .ZN(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4628_ (.A1(_3924_),
    .A2(_4013_),
    .A3(_4208_),
    .A4(_4125_),
    .Z(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4629_ (.A1(_4202_),
    .A2(_4209_),
    .ZN(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4630_ (.A1(_4187_),
    .A2(_4199_),
    .A3(_4210_),
    .ZN(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4631_ (.I(_4211_),
    .Z(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4632_ (.A1(\as2650.r123[1][0] ),
    .A2(_4212_),
    .ZN(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4633_ (.I(_4063_),
    .Z(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4634_ (.I(_4214_),
    .Z(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4635_ (.I(_4215_),
    .Z(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4636_ (.I(_4199_),
    .Z(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4637_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(_3887_),
    .Z(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4638_ (.I(_4218_),
    .Z(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4639_ (.I(_4219_),
    .Z(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4640_ (.I(_4220_),
    .Z(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4641_ (.I(_4221_),
    .Z(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4642_ (.I(_4222_),
    .Z(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4643_ (.A1(_4216_),
    .A2(_4217_),
    .A3(_4223_),
    .ZN(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4644_ (.A1(_4035_),
    .A2(_4185_),
    .B(_4213_),
    .C(_4224_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4645_ (.I(_4035_),
    .Z(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4646_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_3977_),
    .ZN(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4647_ (.A1(_4134_),
    .A2(_4135_),
    .A3(_4226_),
    .Z(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4648_ (.A1(_4047_),
    .A2(_4053_),
    .A3(_4083_),
    .A4(_4089_),
    .Z(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4649_ (.I(_4228_),
    .Z(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4650_ (.A1(_4047_),
    .A2(_4053_),
    .B1(_4083_),
    .B2(_4089_),
    .ZN(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4651_ (.I(_4230_),
    .Z(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4652_ (.A1(_4127_),
    .A2(_4227_),
    .A3(_4229_),
    .A4(_4231_),
    .Z(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4653_ (.I(_4127_),
    .Z(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4654_ (.I(_4228_),
    .Z(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4655_ (.A1(_4233_),
    .A2(_4227_),
    .B1(_4234_),
    .B2(_4231_),
    .ZN(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4656_ (.A1(_4232_),
    .A2(_4235_),
    .ZN(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4657_ (.I(_3924_),
    .Z(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4658_ (.A1(_4228_),
    .A2(_4230_),
    .ZN(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4659_ (.I(_4057_),
    .Z(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4660_ (.A1(_3918_),
    .A2(_4056_),
    .ZN(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4661_ (.A1(_4055_),
    .A2(_4239_),
    .B(_4240_),
    .ZN(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4662_ (.A1(_4238_),
    .A2(_4241_),
    .Z(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4663_ (.A1(_4238_),
    .A2(_4241_),
    .ZN(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4664_ (.A1(_4242_),
    .A2(_4243_),
    .ZN(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4665_ (.I(_4086_),
    .Z(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4666_ (.I(_4245_),
    .Z(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4667_ (.I(_3954_),
    .Z(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4668_ (.A1(_4246_),
    .A2(_4247_),
    .ZN(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4669_ (.A1(_4237_),
    .A2(_4248_),
    .ZN(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4670_ (.I(_4093_),
    .Z(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4671_ (.I(_4075_),
    .Z(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4672_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_4081_),
    .Z(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4673_ (.A1(_4080_),
    .A2(_4252_),
    .ZN(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4674_ (.I(\as2650.r0[2] ),
    .Z(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4675_ (.I(_4254_),
    .Z(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4676_ (.I(_4255_),
    .Z(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4677_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123[0][2] ),
    .I2(\as2650.r123_2[1][2] ),
    .I3(\as2650.r123_2[0][2] ),
    .S0(_3891_),
    .S1(_4045_),
    .Z(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4678_ (.A1(_4256_),
    .A2(_3894_),
    .B1(_4087_),
    .B2(_4257_),
    .ZN(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4679_ (.A1(_4253_),
    .A2(_4258_),
    .ZN(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4680_ (.I(_4259_),
    .Z(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4681_ (.I(_4260_),
    .Z(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4682_ (.I(_4091_),
    .Z(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4683_ (.A1(_3942_),
    .A2(_3989_),
    .ZN(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4684_ (.I(_4263_),
    .Z(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4685_ (.A1(_4134_),
    .A2(_4135_),
    .B(_4018_),
    .ZN(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4686_ (.A1(_4055_),
    .A2(_4264_),
    .B(_4265_),
    .ZN(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4687_ (.A1(_4262_),
    .A2(_4266_),
    .Z(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4688_ (.I(net6),
    .Z(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4689_ (.I(_4268_),
    .Z(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4690_ (.I(_4269_),
    .Z(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4691_ (.I(_4270_),
    .Z(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4692_ (.I(_4271_),
    .Z(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4693_ (.A1(_4272_),
    .A2(_3967_),
    .ZN(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4694_ (.A1(_4072_),
    .A2(_4267_),
    .B(_4273_),
    .C(_4079_),
    .ZN(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4695_ (.A1(_4032_),
    .A2(_4261_),
    .B(_4274_),
    .C(_4111_),
    .ZN(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4696_ (.A1(_4250_),
    .A2(_4251_),
    .B(_4275_),
    .C(_4067_),
    .ZN(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4697_ (.I(_4125_),
    .Z(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4698_ (.A1(_4237_),
    .A2(_4244_),
    .B1(_4249_),
    .B2(_4276_),
    .C(_4277_),
    .ZN(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4699_ (.I(_3988_),
    .Z(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4700_ (.I(_3990_),
    .Z(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4701_ (.A1(_3926_),
    .A2(_4279_),
    .A3(_4280_),
    .A4(_3992_),
    .ZN(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4702_ (.I(_4281_),
    .Z(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4703_ (.A1(_4126_),
    .A2(_4236_),
    .B(_4278_),
    .C(_4282_),
    .ZN(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4704_ (.A1(_4143_),
    .A2(_4145_),
    .ZN(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4705_ (.I(\as2650.holding_reg[1] ),
    .Z(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4706_ (.A1(_4285_),
    .A2(_4188_),
    .ZN(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4707_ (.A1(_4165_),
    .A2(_4084_),
    .A3(_4090_),
    .Z(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4708_ (.A1(_4286_),
    .A2(_4287_),
    .Z(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4709_ (.I(_4288_),
    .Z(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4710_ (.A1(_4284_),
    .A2(_4289_),
    .ZN(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4711_ (.I(_4016_),
    .Z(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4712_ (.A1(_4291_),
    .A2(_4172_),
    .ZN(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4713_ (.I(\as2650.holding_reg[1] ),
    .ZN(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4714_ (.A1(_4084_),
    .A2(_4090_),
    .B(_4293_),
    .ZN(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4715_ (.A1(_4137_),
    .A2(_4141_),
    .B(_4109_),
    .ZN(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4716_ (.A1(_4084_),
    .A2(_4090_),
    .Z(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4717_ (.A1(_4293_),
    .A2(_4296_),
    .Z(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4718_ (.A1(_4167_),
    .A2(_4168_),
    .B(_4152_),
    .ZN(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4719_ (.A1(_4295_),
    .A2(_4297_),
    .A3(_4298_),
    .Z(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4720_ (.A1(_4295_),
    .A2(_4298_),
    .B(_4297_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4721_ (.A1(_4291_),
    .A2(_4175_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4722_ (.A1(_4299_),
    .A2(_0284_),
    .B(_0285_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4723_ (.A1(_4192_),
    .A2(_4171_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4724_ (.A1(_4138_),
    .A2(_4139_),
    .A3(_4140_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4725_ (.A1(_4162_),
    .A2(_0288_),
    .B(_4137_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4726_ (.A1(_4297_),
    .A2(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4727_ (.A1(_3940_),
    .A2(_4092_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4728_ (.A1(_4285_),
    .A2(_4190_),
    .B(_4156_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4729_ (.A1(_4160_),
    .A2(_0290_),
    .B1(_0291_),
    .B2(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4730_ (.A1(_0286_),
    .A2(_0287_),
    .A3(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4731_ (.I(_4296_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4732_ (.A1(_4293_),
    .A2(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4733_ (.A1(_4291_),
    .A2(_0296_),
    .B(_4171_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4734_ (.A1(_0294_),
    .A2(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4735_ (.A1(_4292_),
    .A2(_4294_),
    .B(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4736_ (.A1(_4290_),
    .A2(_0299_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4737_ (.I(_0300_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4738_ (.A1(_4039_),
    .A2(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4739_ (.A1(_4283_),
    .A2(_0302_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4740_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123_2[0][1] ),
    .S(_3886_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4741_ (.I(_0304_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4742_ (.I(_0305_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4743_ (.I(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4744_ (.I(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4745_ (.A1(_4245_),
    .A2(_4063_),
    .A3(_4221_),
    .A4(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4746_ (.I(_4246_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4747_ (.A1(_0310_),
    .A2(_4223_),
    .B1(_0308_),
    .B2(_4215_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4748_ (.I(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4749_ (.A1(_0309_),
    .A2(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4750_ (.I(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4751_ (.A1(\as2650.r123[1][1] ),
    .A2(_4212_),
    .B1(_0314_),
    .B2(_4217_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4752_ (.A1(_4225_),
    .A2(_0303_),
    .B(_0315_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4753_ (.I(_4281_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4754_ (.I(_4284_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4755_ (.I(_4253_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4756_ (.I(_4258_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4757_ (.I(\as2650.holding_reg[2] ),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4758_ (.A1(_0318_),
    .A2(_0319_),
    .B(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4759_ (.A1(_0320_),
    .A2(_0318_),
    .A3(_0319_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4760_ (.A1(_0321_),
    .A2(_0322_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4761_ (.I(_0323_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4762_ (.I(_4160_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4763_ (.A1(_4285_),
    .A2(_4262_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4764_ (.A1(_4285_),
    .A2(_4262_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4765_ (.A1(_0326_),
    .A2(_0289_),
    .B(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4766_ (.A1(_0324_),
    .A2(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4767_ (.A1(_0325_),
    .A2(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4768_ (.I(_0285_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4769_ (.A1(_4288_),
    .A2(_4294_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4770_ (.A1(_0284_),
    .A2(_0332_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4771_ (.A1(_0324_),
    .A2(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4772_ (.I(_4190_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4773_ (.I(_0335_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4774_ (.A1(_0318_),
    .A2(_0319_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4775_ (.I(_0337_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4776_ (.A1(\as2650.holding_reg[2] ),
    .A2(_0335_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4777_ (.A1(_0336_),
    .A2(_0338_),
    .B(_0339_),
    .C(_4176_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4778_ (.A1(_0287_),
    .A2(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4779_ (.A1(_0331_),
    .A2(_0334_),
    .B(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4780_ (.A1(_4154_),
    .A2(_0322_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4781_ (.I(_4172_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4782_ (.A1(_0330_),
    .A2(_0342_),
    .B1(_0343_),
    .B2(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4783_ (.I(_0321_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4784_ (.A1(_4292_),
    .A2(_0346_),
    .B(_4284_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4785_ (.A1(_0317_),
    .A2(_0324_),
    .B1(_0345_),
    .B2(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4786_ (.I(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4787_ (.I(_0295_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4788_ (.I(net7),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4789_ (.I(_0351_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4790_ (.I(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4791_ (.I(_4071_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4792_ (.I(_4073_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4793_ (.A1(_4092_),
    .A2(_4265_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4794_ (.A1(_4264_),
    .A2(_4234_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4795_ (.A1(_0356_),
    .A2(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4796_ (.A1(_0338_),
    .A2(_0358_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4797_ (.A1(_0354_),
    .A2(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4798_ (.A1(_0353_),
    .A2(_0354_),
    .B(_0355_),
    .C(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4799_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_3888_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4800_ (.A1(_4080_),
    .A2(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4801_ (.I(\as2650.r0[3] ),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4802_ (.I(_0364_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4803_ (.I(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4804_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123[0][3] ),
    .I2(\as2650.r123_2[1][3] ),
    .I3(\as2650.r123_2[0][3] ),
    .S0(_3882_),
    .S1(_4081_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4805_ (.A1(_0366_),
    .A2(_3894_),
    .B1(_4087_),
    .B2(_0367_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4806_ (.A1(_0363_),
    .A2(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4807_ (.I(_0369_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4808_ (.A1(_4032_),
    .A2(_0370_),
    .B(_4111_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4809_ (.A1(_4250_),
    .A2(_0350_),
    .B1(_0361_),
    .B2(_0371_),
    .C(_4067_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4810_ (.I(_4256_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4811_ (.I(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4812_ (.A1(_0374_),
    .A2(_4067_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4813_ (.A1(_4237_),
    .A2(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4814_ (.I(_4240_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4815_ (.I(_4259_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4816_ (.A1(_0378_),
    .A2(_4229_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4817_ (.A1(_0378_),
    .A2(_4231_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4818_ (.A1(_4058_),
    .A2(_3919_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4819_ (.I(_4060_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4820_ (.I(_0337_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4821_ (.A1(_0382_),
    .A2(_0383_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4822_ (.A1(_0377_),
    .A2(_0379_),
    .B1(_0380_),
    .B2(_0381_),
    .C(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4823_ (.I(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4824_ (.A1(_4114_),
    .A2(_0386_),
    .B(_4116_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4825_ (.A1(_0372_),
    .A2(_0376_),
    .B(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4826_ (.A1(_4226_),
    .A2(_0379_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4827_ (.A1(_3976_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4828_ (.A1(_4129_),
    .A2(_0383_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4829_ (.A1(_0390_),
    .A2(_0380_),
    .B(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4830_ (.A1(_0389_),
    .A2(_0392_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4831_ (.A1(_4116_),
    .A2(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4832_ (.A1(_4281_),
    .A2(_0388_),
    .A3(_0394_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4833_ (.A1(_0316_),
    .A2(_0349_),
    .B(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4834_ (.A1(_0373_),
    .A2(_4220_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4835_ (.A1(_4245_),
    .A2(_0307_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4836_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123_2[0][2] ),
    .S(\as2650.psl[4] ),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4837_ (.I(_0399_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4838_ (.I(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4839_ (.A1(_4049_),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4840_ (.I(_0401_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4841_ (.A1(_4085_),
    .A2(_4049_),
    .A3(_0305_),
    .A4(_0403_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4842_ (.A1(_0398_),
    .A2(_0402_),
    .B(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4843_ (.A1(_0397_),
    .A2(_0405_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4844_ (.A1(_0309_),
    .A2(_0406_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4845_ (.I(_4199_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4846_ (.A1(\as2650.r123[1][2] ),
    .A2(_4212_),
    .B1(_0407_),
    .B2(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4847_ (.A1(_4225_),
    .A2(_0396_),
    .B(_0409_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4848_ (.I(_0366_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4849_ (.I(_3888_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4850_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4851_ (.A1(_4099_),
    .A2(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4852_ (.I(\as2650.r0[4] ),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4853_ (.I(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4854_ (.I(_0415_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4855_ (.I(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4856_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123[0][4] ),
    .I2(\as2650.r123_2[1][4] ),
    .I3(\as2650.r123_2[0][4] ),
    .S0(_3882_),
    .S1(_3888_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4857_ (.A1(_0417_),
    .A2(_3895_),
    .B1(_4103_),
    .B2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4858_ (.A1(_0413_),
    .A2(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4859_ (.I(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4860_ (.I(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4861_ (.I(net8),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4862_ (.I(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4863_ (.I(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4864_ (.I(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4865_ (.I(_0426_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4866_ (.A1(_0363_),
    .A2(_0368_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4867_ (.I(_0428_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4868_ (.A1(_4262_),
    .A2(_4260_),
    .A3(_4265_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4869_ (.A1(_0337_),
    .A2(_4263_),
    .A3(_4229_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4870_ (.A1(_0430_),
    .A2(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4871_ (.A1(_0429_),
    .A2(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4872_ (.A1(_4072_),
    .A2(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4873_ (.A1(_0427_),
    .A2(_0354_),
    .B(_0355_),
    .C(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4874_ (.I(_4014_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4875_ (.I(_0436_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4876_ (.I(_0437_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4877_ (.I(_4020_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4878_ (.A1(_0438_),
    .A2(_3898_),
    .A3(_3965_),
    .A4(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4879_ (.A1(_0355_),
    .A2(_0422_),
    .B(_0435_),
    .C(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4880_ (.I(_0338_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4881_ (.A1(_4250_),
    .A2(_0442_),
    .B(_4247_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4882_ (.A1(_0410_),
    .A2(_4066_),
    .B1(_0441_),
    .B2(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4883_ (.A1(_0318_),
    .A2(_0319_),
    .A3(_0363_),
    .A4(_0368_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4884_ (.A1(_4229_),
    .A2(_0445_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4885_ (.I(_0428_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4886_ (.A1(_0383_),
    .A2(_4234_),
    .B(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4887_ (.A1(_0446_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4888_ (.A1(_0378_),
    .A2(_4231_),
    .A3(_0369_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4889_ (.A1(_4075_),
    .A2(_0295_),
    .A3(_0383_),
    .B(_0447_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4890_ (.A1(_0450_),
    .A2(_0451_),
    .B(_0381_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4891_ (.A1(_0382_),
    .A2(_0429_),
    .B1(_0449_),
    .B2(_4059_),
    .C(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4892_ (.I(_0453_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4893_ (.A1(_4043_),
    .A2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4894_ (.I(_4125_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4895_ (.A1(_4043_),
    .A2(_0444_),
    .B(_0455_),
    .C(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4896_ (.A1(_0450_),
    .A2(_0451_),
    .B(_0390_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4897_ (.A1(_4129_),
    .A2(_0429_),
    .B1(_0449_),
    .B2(_4128_),
    .C(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4898_ (.I(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4899_ (.A1(_4116_),
    .A2(_0460_),
    .B(_4038_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4900_ (.I(\as2650.holding_reg[3] ),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4901_ (.A1(_0462_),
    .A2(_3937_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4902_ (.I(\as2650.holding_reg[3] ),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4903_ (.A1(_0363_),
    .A2(_0368_),
    .B(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4904_ (.A1(_3937_),
    .A2(_0428_),
    .B(_0463_),
    .C(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4905_ (.A1(_0462_),
    .A2(_4188_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4906_ (.A1(_4188_),
    .A2(_0428_),
    .B(_0465_),
    .C(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4907_ (.A1(_0466_),
    .A2(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4908_ (.I(_0469_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4909_ (.I(_4189_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4910_ (.A1(_0471_),
    .A2(_0447_),
    .B(_0467_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4911_ (.I(_4176_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4912_ (.A1(_0464_),
    .A2(_4189_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4913_ (.A1(_0471_),
    .A2(_0369_),
    .B(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4914_ (.A1(\as2650.holding_reg[2] ),
    .A2(_3938_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4915_ (.A1(_3938_),
    .A2(_0337_),
    .B(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4916_ (.I(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4917_ (.A1(_0284_),
    .A2(_0332_),
    .B(_0324_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4918_ (.A1(_0346_),
    .A2(_0478_),
    .B(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4919_ (.A1(_0470_),
    .A2(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4920_ (.A1(_4291_),
    .A2(_4156_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4921_ (.A1(_0320_),
    .A2(_0338_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4922_ (.A1(_0483_),
    .A2(_0328_),
    .B(_0346_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4923_ (.A1(_0470_),
    .A2(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4924_ (.A1(_0482_),
    .A2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4925_ (.A1(_0473_),
    .A2(_0475_),
    .B1(_0481_),
    .B2(_0331_),
    .C(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4926_ (.A1(_4172_),
    .A2(_0472_),
    .B(_0487_),
    .C(_4148_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4927_ (.I(_4292_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4928_ (.A1(_0489_),
    .A2(_0465_),
    .B(_4284_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4929_ (.A1(_0317_),
    .A2(_0470_),
    .B1(_0488_),
    .B2(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4930_ (.I(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4931_ (.A1(_0457_),
    .A2(_0461_),
    .B1(_0492_),
    .B2(_4039_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4932_ (.A1(_3896_),
    .A2(_3941_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4933_ (.A1(_4143_),
    .A2(_0494_),
    .A3(_4194_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4934_ (.A1(_4023_),
    .A2(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4935_ (.I(\as2650.r0[1] ),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4936_ (.I(_0400_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4937_ (.A1(_0497_),
    .A2(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4938_ (.A1(_0373_),
    .A2(_0307_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4939_ (.I(_0403_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4940_ (.A1(_4256_),
    .A2(_4086_),
    .A3(_0306_),
    .A4(_0501_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4941_ (.A1(_0499_),
    .A2(_0500_),
    .B(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4942_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123_2[0][3] ),
    .S(_3887_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4943_ (.I(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4944_ (.A1(_4050_),
    .A2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4945_ (.A1(_0366_),
    .A2(_4219_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4946_ (.A1(_0404_),
    .A2(_0506_),
    .A3(_0507_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4947_ (.A1(_0503_),
    .A2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4948_ (.A1(_0373_),
    .A2(_4222_),
    .A3(_0405_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4949_ (.A1(_0309_),
    .A2(_0406_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4950_ (.A1(_0510_),
    .A2(_0511_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4951_ (.A1(_0509_),
    .A2(_0512_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4952_ (.A1(_0496_),
    .A2(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4953_ (.A1(\as2650.r123[1][3] ),
    .A2(_4212_),
    .B(_0514_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4954_ (.A1(_4225_),
    .A2(_0493_),
    .B(_0515_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4955_ (.I(\as2650.holding_reg[4] ),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4956_ (.A1(_0516_),
    .A2(_4166_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4957_ (.A1(_4189_),
    .A2(_0420_),
    .B(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4958_ (.I(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4959_ (.A1(_4166_),
    .A2(_0420_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4960_ (.A1(\as2650.holding_reg[4] ),
    .A2(_4166_),
    .B(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4961_ (.A1(_0519_),
    .A2(_0521_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4962_ (.I(_0429_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4963_ (.A1(_0464_),
    .A2(_0523_),
    .B1(_0470_),
    .B2(_0484_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4964_ (.A1(_0522_),
    .A2(_0524_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4965_ (.A1(_0325_),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4966_ (.A1(_0518_),
    .A2(_0521_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4967_ (.A1(_4286_),
    .A2(_4287_),
    .A3(_4294_),
    .B1(_0346_),
    .B2(_0322_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4968_ (.A1(_0466_),
    .A2(_0468_),
    .A3(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4969_ (.A1(_4289_),
    .A2(_0296_),
    .B(_4298_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4970_ (.A1(_0322_),
    .A2(_0468_),
    .A3(_0477_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4971_ (.A1(_0475_),
    .A2(_0472_),
    .B1(_0529_),
    .B2(_0530_),
    .C(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4972_ (.A1(_0284_),
    .A2(_0332_),
    .B(_0469_),
    .C(_0323_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4973_ (.A1(_0532_),
    .A2(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4974_ (.A1(_0527_),
    .A2(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4975_ (.A1(_4156_),
    .A2(_0519_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4976_ (.A1(_0331_),
    .A2(_0535_),
    .B(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4977_ (.I(_4154_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4978_ (.I(_0521_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4979_ (.A1(_0538_),
    .A2(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4980_ (.A1(_0526_),
    .A2(_0537_),
    .B1(_0540_),
    .B2(_0344_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4981_ (.A1(_0413_),
    .A2(_0419_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4982_ (.I(_0542_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4983_ (.I(_0543_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4984_ (.A1(_0516_),
    .A2(_0544_),
    .B(_0489_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4985_ (.A1(_4147_),
    .A2(_0527_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4986_ (.A1(_4147_),
    .A2(_0541_),
    .A3(_0545_),
    .B(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4987_ (.I(_0547_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4988_ (.I(_4129_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4989_ (.A1(_0543_),
    .A2(_0450_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4990_ (.A1(_4228_),
    .A2(_0420_),
    .A3(_0445_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4991_ (.I(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4992_ (.A1(_4234_),
    .A2(_0445_),
    .B(_0421_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4993_ (.A1(_4226_),
    .A2(_0552_),
    .A3(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4994_ (.A1(_0549_),
    .A2(_0421_),
    .B1(_0550_),
    .B2(_4233_),
    .C(_0554_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4995_ (.I(_0555_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4996_ (.I(_0417_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4997_ (.I(net9),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4998_ (.I(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4999_ (.I(_0559_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5000_ (.I(_0560_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5001_ (.I(_4071_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5002_ (.I0(_0430_),
    .I1(_0431_),
    .S(_0447_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5003_ (.A1(_0543_),
    .A2(_0563_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5004_ (.A1(_3967_),
    .A2(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5005_ (.A1(_0561_),
    .A2(_0562_),
    .B(_4074_),
    .C(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5006_ (.I(\as2650.r123_2[1][5] ),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5007_ (.A1(_3889_),
    .A2(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5008_ (.I(_3892_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5009_ (.A1(_0411_),
    .A2(\as2650.r123[1][5] ),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5010_ (.A1(_3883_),
    .A2(_0569_),
    .A3(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5011_ (.I0(\as2650.r123[0][5] ),
    .I1(\as2650.r123_2[0][5] ),
    .S(_3886_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5012_ (.I(_0572_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5013_ (.I(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5014_ (.A1(_3884_),
    .A2(_3892_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5015_ (.A1(_0568_),
    .A2(_0571_),
    .B1(_0574_),
    .B2(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5016_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_0411_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5017_ (.A1(_4099_),
    .A2(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5018_ (.I(\as2650.r0[5] ),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5019_ (.I(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5020_ (.I(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5021_ (.A1(_0581_),
    .A2(_3895_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5022_ (.A1(_0576_),
    .A2(_0578_),
    .A3(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5023_ (.I(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5024_ (.I(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5025_ (.I(_0585_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5026_ (.A1(_4079_),
    .A2(_0586_),
    .B(_4093_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5027_ (.A1(_4022_),
    .A2(_0523_),
    .B1(_0566_),
    .B2(_0587_),
    .C(_4065_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5028_ (.A1(_0557_),
    .A2(_4247_),
    .B(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5029_ (.A1(_0377_),
    .A2(_0552_),
    .A3(_0553_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5030_ (.A1(_0381_),
    .A2(_0377_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5031_ (.A1(_0591_),
    .A2(_0543_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5032_ (.A1(_4239_),
    .A2(_0550_),
    .B(_0590_),
    .C(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5033_ (.I(_0593_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5034_ (.A1(_4042_),
    .A2(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5035_ (.A1(_4114_),
    .A2(_0589_),
    .B(_0595_),
    .C(_4277_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5036_ (.A1(_0456_),
    .A2(_0556_),
    .B(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5037_ (.A1(_4282_),
    .A2(_0597_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5038_ (.A1(_0316_),
    .A2(_0548_),
    .B(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5039_ (.I(_4211_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5040_ (.A1(_0511_),
    .A2(_0509_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5041_ (.A1(_0510_),
    .A2(_0509_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5042_ (.A1(_0503_),
    .A2(_0508_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5043_ (.I(_0506_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5044_ (.A1(_4245_),
    .A2(_4063_),
    .A3(_0307_),
    .A4(_0501_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5045_ (.A1(_0605_),
    .A2(_0507_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5046_ (.A1(_0605_),
    .A2(_0507_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5047_ (.A1(_0604_),
    .A2(_0606_),
    .B(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5048_ (.A1(_4255_),
    .A2(_0498_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5049_ (.A1(_0365_),
    .A2(_0305_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5050_ (.I0(\as2650.r123[0][4] ),
    .I1(\as2650.r123_2[0][4] ),
    .S(\as2650.psl[4] ),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5051_ (.I(_0611_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5052_ (.I(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5053_ (.I(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5054_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5055_ (.A1(_4050_),
    .A2(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5056_ (.A1(_0609_),
    .A2(_0610_),
    .A3(_0616_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5057_ (.A1(_4256_),
    .A2(_4086_),
    .A3(_0306_),
    .A4(_0403_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5058_ (.A1(_4085_),
    .A2(_0505_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5059_ (.A1(_0416_),
    .A2(_4220_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5060_ (.A1(_0618_),
    .A2(_0619_),
    .A3(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5061_ (.A1(_0617_),
    .A2(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5062_ (.A1(_0603_),
    .A2(_0608_),
    .A3(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5063_ (.A1(_0601_),
    .A2(_0602_),
    .A3(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5064_ (.A1(\as2650.r123[1][4] ),
    .A2(_0600_),
    .B1(_0624_),
    .B2(_0408_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5065_ (.A1(_4225_),
    .A2(_0599_),
    .B(_0625_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5066_ (.I(_0317_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5067_ (.I(\as2650.holding_reg[5] ),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5068_ (.A1(_0627_),
    .A2(_0585_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5069_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0584_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5070_ (.A1(_0628_),
    .A2(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5071_ (.A1(_0519_),
    .A2(_0521_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5072_ (.A1(_0532_),
    .A2(_0533_),
    .B(_0527_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5073_ (.A1(_0631_),
    .A2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5074_ (.A1(_0630_),
    .A2(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5075_ (.A1(_0516_),
    .A2(_0544_),
    .B1(_0527_),
    .B2(_0524_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5076_ (.A1(_0630_),
    .A2(_0635_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5077_ (.A1(_0576_),
    .A2(_0578_),
    .A3(_0582_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5078_ (.I(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5079_ (.I(_0638_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5080_ (.A1(_0627_),
    .A2(_0336_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5081_ (.A1(_0336_),
    .A2(_0639_),
    .B(_0640_),
    .C(_4176_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5082_ (.A1(_0482_),
    .A2(_0636_),
    .B(_0641_),
    .C(_0287_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5083_ (.A1(_0331_),
    .A2(_0634_),
    .B(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5084_ (.A1(_0344_),
    .A2(_0629_),
    .B(_0643_),
    .C(_4148_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5085_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0584_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5086_ (.A1(_0489_),
    .A2(_0645_),
    .B(_0317_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5087_ (.A1(_0626_),
    .A2(_0630_),
    .B1(_0644_),
    .B2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5088_ (.I(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5089_ (.A1(_0552_),
    .A2(_0638_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5090_ (.A1(_0378_),
    .A2(_4230_),
    .A3(_0369_),
    .A4(_0542_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5091_ (.A1(_0650_),
    .A2(_0583_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5092_ (.A1(_0390_),
    .A2(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5093_ (.A1(_0549_),
    .A2(_0638_),
    .B1(_0649_),
    .B2(_4128_),
    .C(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5094_ (.I(_0653_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5095_ (.I(_0581_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5096_ (.I(net1),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5097_ (.I(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5098_ (.I(_0657_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5099_ (.A1(_3899_),
    .A2(_3945_),
    .A3(_3947_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5100_ (.A1(_3944_),
    .A2(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5101_ (.A1(_4264_),
    .A2(_0552_),
    .B1(_0650_),
    .B2(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5102_ (.A1(_0585_),
    .A2(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5103_ (.A1(_4071_),
    .A2(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5104_ (.A1(_0658_),
    .A2(_0562_),
    .B(_4073_),
    .C(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5105_ (.I(\as2650.r0[6] ),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5106_ (.I(_0665_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5107_ (.I(_0666_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5108_ (.A1(_0667_),
    .A2(_3895_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5109_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_0411_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5110_ (.A1(_4099_),
    .A2(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5111_ (.I0(\as2650.r123[1][6] ),
    .I1(\as2650.r123[0][6] ),
    .I2(\as2650.r123_2[1][6] ),
    .I3(\as2650.r123_2[0][6] ),
    .S0(_3883_),
    .S1(_3889_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5112_ (.A1(_4103_),
    .A2(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5113_ (.A1(_0668_),
    .A2(_0670_),
    .A3(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5114_ (.I(_0673_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5115_ (.I(_0674_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5116_ (.I(_0675_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5117_ (.A1(_4079_),
    .A2(_0676_),
    .B(_4093_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5118_ (.A1(_4022_),
    .A2(_0422_),
    .B1(_0664_),
    .B2(_0677_),
    .C(_3954_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5119_ (.A1(_0655_),
    .A2(_4247_),
    .B(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5120_ (.A1(_0381_),
    .A2(_0651_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5121_ (.A1(_0382_),
    .A2(_0639_),
    .B1(_0649_),
    .B2(_4059_),
    .C(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5122_ (.I(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5123_ (.A1(_4042_),
    .A2(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5124_ (.A1(_4042_),
    .A2(_0679_),
    .B(_0683_),
    .C(_4277_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5125_ (.A1(_0456_),
    .A2(_0654_),
    .B(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5126_ (.A1(_4282_),
    .A2(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5127_ (.A1(_0316_),
    .A2(_0648_),
    .B(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5128_ (.A1(_0602_),
    .A2(_0623_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5129_ (.A1(_0602_),
    .A2(_0623_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5130_ (.A1(_0601_),
    .A2(_0688_),
    .B(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5131_ (.A1(_0603_),
    .A2(_0622_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5132_ (.A1(_0603_),
    .A2(_0622_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5133_ (.A1(_0608_),
    .A2(_0691_),
    .B(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5134_ (.A1(_0617_),
    .A2(_0621_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5135_ (.A1(_0618_),
    .A2(_0620_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5136_ (.A1(_0417_),
    .A2(_4220_),
    .A3(_0502_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5137_ (.A1(_0619_),
    .A2(_0695_),
    .B(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5138_ (.A1(_4049_),
    .A2(_0573_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5139_ (.A1(_0414_),
    .A2(_0304_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5140_ (.A1(\as2650.r0[1] ),
    .A2(_0612_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5141_ (.A1(_0365_),
    .A2(_0401_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5142_ (.A1(_0699_),
    .A2(_0700_),
    .A3(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5143_ (.A1(_0698_),
    .A2(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5144_ (.A1(_4255_),
    .A2(_0505_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5145_ (.A1(\as2650.r0[2] ),
    .A2(_0611_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5146_ (.A1(_4255_),
    .A2(_0401_),
    .B1(_0613_),
    .B2(_4048_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5147_ (.A1(_0402_),
    .A2(_0705_),
    .B1(_0706_),
    .B2(_0610_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5148_ (.A1(_0579_),
    .A2(_4219_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5149_ (.A1(_0704_),
    .A2(_0707_),
    .A3(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5150_ (.A1(_0703_),
    .A2(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5151_ (.A1(_0694_),
    .A2(_0697_),
    .A3(_0710_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5152_ (.A1(_0690_),
    .A2(_0693_),
    .A3(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5153_ (.A1(\as2650.r123[1][5] ),
    .A2(_0600_),
    .B1(_0712_),
    .B2(_0408_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5154_ (.A1(_4035_),
    .A2(_0687_),
    .B(_0713_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5155_ (.A1(_0668_),
    .A2(_0670_),
    .A3(_0672_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5156_ (.I(_0714_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5157_ (.A1(_0650_),
    .A2(_0584_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5158_ (.A1(_0674_),
    .A2(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5159_ (.A1(_0551_),
    .A2(_0637_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5160_ (.A1(_0674_),
    .A2(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5161_ (.A1(_4226_),
    .A2(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5162_ (.A1(_0549_),
    .A2(_0715_),
    .B1(_0717_),
    .B2(_4233_),
    .C(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5163_ (.I(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5164_ (.A1(_0456_),
    .A2(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5165_ (.A1(_0377_),
    .A2(_0719_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5166_ (.A1(_0382_),
    .A2(_0715_),
    .B1(_0717_),
    .B2(_4239_),
    .C(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5167_ (.I(_0725_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5168_ (.I(net2),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5169_ (.I(_0727_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5170_ (.I(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5171_ (.I(_0729_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5172_ (.A1(_4264_),
    .A2(_0551_),
    .A3(_0637_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5173_ (.A1(_4018_),
    .A2(_0716_),
    .B(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5174_ (.A1(_0675_),
    .A2(_0732_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5175_ (.A1(_0562_),
    .A2(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5176_ (.A1(_0730_),
    .A2(_4072_),
    .B(_4074_),
    .C(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5177_ (.A1(_4098_),
    .A2(_4102_),
    .A3(_4105_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5178_ (.I(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5179_ (.I(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5180_ (.A1(_4032_),
    .A2(_0738_),
    .B(_4022_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5181_ (.A1(_4111_),
    .A2(_0586_),
    .B1(_0735_),
    .B2(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5182_ (.I(_0667_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5183_ (.A1(_0741_),
    .A2(_4065_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5184_ (.A1(_4066_),
    .A2(_0740_),
    .B(_0742_),
    .C(_3924_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5185_ (.A1(_4237_),
    .A2(_0726_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5186_ (.A1(_4126_),
    .A2(_0744_),
    .B(_4038_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5187_ (.A1(\as2650.holding_reg[6] ),
    .A2(_3939_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5188_ (.A1(_3939_),
    .A2(_0714_),
    .B(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5189_ (.A1(_3939_),
    .A2(_0714_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5190_ (.A1(\as2650.holding_reg[6] ),
    .A2(_3940_),
    .B(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5191_ (.A1(_0747_),
    .A2(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5192_ (.A1(_0747_),
    .A2(_0749_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5193_ (.A1(_0750_),
    .A2(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5194_ (.I(\as2650.holding_reg[6] ),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5195_ (.A1(_0750_),
    .A2(_0751_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5196_ (.A1(_0627_),
    .A2(_0585_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5197_ (.A1(_0755_),
    .A2(_0635_),
    .B(_0628_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5198_ (.A1(_0754_),
    .A2(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5199_ (.A1(_0471_),
    .A2(_0637_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5200_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0471_),
    .B(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5201_ (.A1(_0645_),
    .A2(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5202_ (.A1(_0629_),
    .A2(_0759_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5203_ (.A1(_0631_),
    .A2(_0632_),
    .A3(_0760_),
    .B(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5204_ (.A1(_0752_),
    .A2(_0762_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5205_ (.A1(_4157_),
    .A2(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5206_ (.A1(_0473_),
    .A2(_0749_),
    .B1(_0757_),
    .B2(_0325_),
    .C(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5207_ (.A1(_0753_),
    .A2(_0287_),
    .A3(_0676_),
    .B1(_0765_),
    .B2(_0344_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5208_ (.A1(_0753_),
    .A2(_0676_),
    .B(_0489_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5209_ (.A1(_0766_),
    .A2(_0767_),
    .B(_0626_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5210_ (.A1(_0626_),
    .A2(_0752_),
    .B(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5211_ (.A1(_4281_),
    .A2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5212_ (.A1(_0723_),
    .A2(_0745_),
    .B(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5213_ (.A1(_0693_),
    .A2(_0711_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5214_ (.A1(_0693_),
    .A2(_0711_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5215_ (.A1(_0690_),
    .A2(_0772_),
    .B(_0773_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5216_ (.A1(_0694_),
    .A2(_0710_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5217_ (.A1(_0694_),
    .A2(_0710_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5218_ (.A1(_0697_),
    .A2(_0775_),
    .B(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5219_ (.A1(_0581_),
    .A2(_4221_),
    .B(_0707_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5220_ (.A1(_0581_),
    .A2(_4221_),
    .A3(_0707_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5221_ (.A1(_0704_),
    .A2(_0778_),
    .B(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5222_ (.A1(_0703_),
    .A2(_0709_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5223_ (.A1(_0698_),
    .A2(_0702_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5224_ (.A1(_4085_),
    .A2(_0573_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5225_ (.I0(\as2650.r123[0][6] ),
    .I1(\as2650.r123_2[0][6] ),
    .S(\as2650.psl[4] ),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5226_ (.I(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5227_ (.I(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5228_ (.A1(_4048_),
    .A2(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5229_ (.I(_0572_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5230_ (.A1(_0497_),
    .A2(_4048_),
    .A3(_0788_),
    .A4(_0785_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5231_ (.A1(_0783_),
    .A2(_0787_),
    .B(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5232_ (.A1(\as2650.r0[5] ),
    .A2(_0304_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5233_ (.A1(_0414_),
    .A2(_0400_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5234_ (.A1(_0705_),
    .A2(_0791_),
    .A3(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5235_ (.A1(_0790_),
    .A2(_0793_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5236_ (.A1(_0365_),
    .A2(_0504_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5237_ (.A1(_0364_),
    .A2(_0611_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5238_ (.A1(_0364_),
    .A2(_0498_),
    .B1(_0612_),
    .B2(_0497_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5239_ (.A1(_0499_),
    .A2(_0796_),
    .B1(_0797_),
    .B2(_0699_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5240_ (.A1(_0665_),
    .A2(_4218_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5241_ (.I(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5242_ (.A1(_0795_),
    .A2(_0798_),
    .A3(_0800_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5243_ (.A1(_0782_),
    .A2(_0794_),
    .A3(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5244_ (.A1(_0781_),
    .A2(_0802_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5245_ (.A1(_0780_),
    .A2(_0803_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5246_ (.A1(_0777_),
    .A2(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5247_ (.A1(_0774_),
    .A2(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5248_ (.A1(\as2650.r123[1][6] ),
    .A2(_0600_),
    .B1(_0806_),
    .B2(_0408_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5249_ (.A1(_4035_),
    .A2(_0771_),
    .B(_0807_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5250_ (.A1(_0777_),
    .A2(_0804_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5251_ (.A1(_0774_),
    .A2(_0805_),
    .B(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5252_ (.A1(_0781_),
    .A2(_0802_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5253_ (.A1(_0780_),
    .A2(_0803_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5254_ (.A1(_0810_),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5255_ (.A1(_0798_),
    .A2(_0800_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5256_ (.A1(_0798_),
    .A2(_0800_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5257_ (.A1(_0795_),
    .A2(_0813_),
    .B(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5258_ (.A1(_0782_),
    .A2(_0794_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5259_ (.A1(_0782_),
    .A2(_0794_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5260_ (.A1(_0816_),
    .A2(_0801_),
    .B(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5261_ (.A1(_0790_),
    .A2(_0793_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5262_ (.A1(\as2650.r0[6] ),
    .A2(_0305_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5263_ (.A1(\as2650.r0[5] ),
    .A2(_0399_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5264_ (.A1(_0796_),
    .A2(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5265_ (.A1(_0820_),
    .A2(_0822_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5266_ (.A1(\as2650.r0[1] ),
    .A2(_0785_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5267_ (.A1(\as2650.r0[2] ),
    .A2(_0572_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5268_ (.I0(\as2650.r123[0][7] ),
    .I1(\as2650.r123_2[0][7] ),
    .S(_3886_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5269_ (.A1(\as2650.r0[0] ),
    .A2(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5270_ (.A1(_0824_),
    .A2(_0825_),
    .A3(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5271_ (.A1(_0789_),
    .A2(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5272_ (.A1(_0819_),
    .A2(_0823_),
    .A3(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5273_ (.I(_0504_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(_0416_),
    .A2(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5275_ (.A1(_0415_),
    .A2(_0613_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5276_ (.A1(_0415_),
    .A2(_0498_),
    .B1(_0613_),
    .B2(_4254_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5277_ (.A1(_0609_),
    .A2(_0833_),
    .B1(_0834_),
    .B2(_0791_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5278_ (.A1(\as2650.r0[7] ),
    .A2(_4219_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5279_ (.A1(_0835_),
    .A2(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5280_ (.A1(_0832_),
    .A2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5281_ (.A1(_0830_),
    .A2(_0838_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5282_ (.A1(_0818_),
    .A2(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5283_ (.A1(_0815_),
    .A2(_0840_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5284_ (.A1(_0812_),
    .A2(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5285_ (.A1(_0809_),
    .A2(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5286_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0737_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5287_ (.I(_0844_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5288_ (.A1(_0753_),
    .A2(_0675_),
    .B1(_0752_),
    .B2(_0756_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5289_ (.A1(_0845_),
    .A2(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5290_ (.A1(_0752_),
    .A2(_0762_),
    .B(_0750_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5291_ (.A1(_0844_),
    .A2(_0848_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5292_ (.I(_0336_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5293_ (.I(_0335_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5294_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5295_ (.A1(_0850_),
    .A2(_0737_),
    .B(_0852_),
    .C(_0473_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5296_ (.A1(_4157_),
    .A2(_0849_),
    .B(_0853_),
    .C(_4027_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5297_ (.A1(_0325_),
    .A2(_0847_),
    .B(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5298_ (.I(\as2650.holding_reg[7] ),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5299_ (.A1(_0856_),
    .A2(_4107_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5300_ (.A1(_0856_),
    .A2(_4107_),
    .B(_0538_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5301_ (.A1(_4027_),
    .A2(_0857_),
    .A3(_0858_),
    .B(_0626_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5302_ (.A1(_4147_),
    .A2(_0845_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5303_ (.A1(_0855_),
    .A2(_0859_),
    .B(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5304_ (.I(_0861_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5305_ (.A1(_0650_),
    .A2(_0583_),
    .A3(_0674_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5306_ (.A1(_4106_),
    .A2(_0863_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5307_ (.A1(_0542_),
    .A2(_0583_),
    .A3(_0673_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5308_ (.A1(_0446_),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5309_ (.A1(_4106_),
    .A2(_0866_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _5310_ (.A1(_0736_),
    .A2(_0549_),
    .B1(_0864_),
    .B2(_4233_),
    .C1(_0867_),
    .C2(_4128_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5311_ (.I(_4097_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5312_ (.I(_0869_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5313_ (.A1(_4139_),
    .A2(_4140_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5314_ (.I(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5315_ (.A1(_4095_),
    .A2(_0872_),
    .B(_4109_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5316_ (.I(net3),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5317_ (.I(_0874_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5318_ (.I(_0875_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5319_ (.A1(_3943_),
    .A2(_3990_),
    .A3(_0866_),
    .B1(_0863_),
    .B2(_4018_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5320_ (.A1(_0736_),
    .A2(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5321_ (.A1(_0562_),
    .A2(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5322_ (.A1(_0876_),
    .A2(_0354_),
    .B(_4074_),
    .C(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5323_ (.A1(_0355_),
    .A2(_0873_),
    .B(_0880_),
    .C(_0440_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5324_ (.A1(_4250_),
    .A2(_0715_),
    .B(_4065_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5325_ (.A1(_0870_),
    .A2(_4066_),
    .B1(_0881_),
    .B2(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5326_ (.A1(_4106_),
    .A2(_0591_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5327_ (.A1(_4239_),
    .A2(_0864_),
    .B1(_0867_),
    .B2(_4059_),
    .C(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5328_ (.I(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5329_ (.A1(_4114_),
    .A2(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5330_ (.A1(_4043_),
    .A2(_0883_),
    .B(_0887_),
    .C(_4277_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5331_ (.A1(_4126_),
    .A2(_0868_),
    .B(_0888_),
    .C(_4282_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5332_ (.A1(_0316_),
    .A2(_0862_),
    .B(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5333_ (.A1(\as2650.r123[1][7] ),
    .A2(_0600_),
    .B1(_0890_),
    .B2(_4210_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5334_ (.A1(_0496_),
    .A2(_0843_),
    .B(_0891_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5335_ (.I(_0569_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5336_ (.A1(_0892_),
    .A2(_4034_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5337_ (.I(_3935_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5338_ (.A1(_4200_),
    .A2(_0569_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5339_ (.A1(_4192_),
    .A2(_4190_),
    .A3(_4193_),
    .A4(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5340_ (.A1(_3944_),
    .A2(_3996_),
    .A3(_4144_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5341_ (.I(_0897_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5342_ (.A1(_4120_),
    .A2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5343_ (.A1(_0494_),
    .A2(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5344_ (.A1(_0896_),
    .A2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5345_ (.I(_0901_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5346_ (.I(_0902_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5347_ (.I(_0903_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5348_ (.A1(_0894_),
    .A2(_0904_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5349_ (.I(_4000_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5350_ (.A1(_0906_),
    .A2(_4209_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5351_ (.I(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5352_ (.A1(_4187_),
    .A2(_0905_),
    .A3(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5353_ (.A1(_4120_),
    .A2(_0897_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5354_ (.I(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5355_ (.A1(_4191_),
    .A2(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5356_ (.I(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5357_ (.A1(_0894_),
    .A2(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5358_ (.I(\as2650.psu[0] ),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5359_ (.I(\as2650.psu[1] ),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5360_ (.A1(_0915_),
    .A2(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5361_ (.I(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5362_ (.I(_0918_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5363_ (.I(_0919_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5364_ (.I(_0917_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5365_ (.I(\as2650.psu[0] ),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5366_ (.I(\as2650.psu[1] ),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5367_ (.A1(_0922_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5368_ (.I(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5369_ (.A1(_0921_),
    .A2(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5370_ (.I(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5371_ (.I(_0915_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5372_ (.I(_0928_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5373_ (.I0(\as2650.stack[1][8] ),
    .I1(\as2650.stack[0][8] ),
    .S(_0929_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5374_ (.A1(\as2650.stack[2][8] ),
    .A2(_0920_),
    .B1(_0927_),
    .B2(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5375_ (.I(\as2650.psu[2] ),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5376_ (.A1(_0932_),
    .A2(_0925_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5377_ (.I(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5378_ (.I(_0923_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5379_ (.A1(_0922_),
    .A2(_0935_),
    .B(\as2650.psu[2] ),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5380_ (.I(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5381_ (.A1(\as2650.stack[3][8] ),
    .A2(_0934_),
    .B(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5382_ (.I(_0921_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5383_ (.I(_0939_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5384_ (.I(_0935_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5385_ (.I(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5386_ (.I(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5387_ (.I(_0922_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5388_ (.I(_0944_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5389_ (.I(_0945_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5390_ (.A1(_0943_),
    .A2(\as2650.stack[5][8] ),
    .B1(\as2650.stack[4][8] ),
    .B2(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5391_ (.A1(_0940_),
    .A2(_0947_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5392_ (.I(\as2650.psu[2] ),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5393_ (.I(_0949_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5394_ (.I(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5395_ (.A1(_0936_),
    .A2(_0933_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5396_ (.I(_0952_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5397_ (.I(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5398_ (.A1(_0951_),
    .A2(\as2650.stack[7][8] ),
    .B1(\as2650.stack[6][8] ),
    .B2(_0940_),
    .C(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5399_ (.A1(_0931_),
    .A2(_0938_),
    .B1(_0948_),
    .B2(_0955_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5400_ (.I(_0913_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5401_ (.A1(_4197_),
    .A2(_0904_),
    .B(_0894_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5402_ (.A1(_4215_),
    .A2(_0914_),
    .B1(_0956_),
    .B2(_0957_),
    .C(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5403_ (.A1(_0909_),
    .A2(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5404_ (.A1(\as2650.r123[0][0] ),
    .A2(_0909_),
    .B(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5405_ (.A1(_4185_),
    .A2(_0893_),
    .B(_0961_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5406_ (.A1(_4186_),
    .A2(_0905_),
    .A3(_0907_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5407_ (.I(_0962_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5408_ (.A1(\as2650.r123[0][1] ),
    .A2(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5409_ (.I(_0310_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5410_ (.I(_0914_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5411_ (.I(_0919_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5412_ (.I(_0945_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5413_ (.A1(_0943_),
    .A2(\as2650.stack[5][9] ),
    .B1(\as2650.stack[4][9] ),
    .B2(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5414_ (.A1(_0967_),
    .A2(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5415_ (.I(_0952_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5416_ (.I(_0971_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5417_ (.I(_0972_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5418_ (.A1(_0951_),
    .A2(\as2650.stack[7][9] ),
    .B1(\as2650.stack[6][9] ),
    .B2(_0920_),
    .C(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5419_ (.A1(_0936_),
    .A2(_0933_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5420_ (.I(_0975_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5421_ (.I(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5422_ (.I(_0916_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5423_ (.I0(\as2650.stack[3][9] ),
    .I1(\as2650.stack[0][9] ),
    .I2(\as2650.stack[1][9] ),
    .I3(\as2650.stack[2][9] ),
    .S0(_0929_),
    .S1(_0978_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5424_ (.A1(_0977_),
    .A2(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5425_ (.A1(_0970_),
    .A2(_0974_),
    .B(_0980_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5426_ (.I(_0957_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5427_ (.I(_0958_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5428_ (.A1(_0965_),
    .A2(_0966_),
    .B1(_0981_),
    .B2(_0982_),
    .C(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5429_ (.A1(_4283_),
    .A2(_0302_),
    .A3(_0908_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5430_ (.A1(_0963_),
    .A2(_0984_),
    .A3(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5431_ (.A1(_0964_),
    .A2(_0986_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5432_ (.I(_0962_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5433_ (.A1(\as2650.r123[0][2] ),
    .A2(_0987_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5434_ (.I(_0908_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5435_ (.I(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5436_ (.I(_0962_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5437_ (.I(_0374_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5438_ (.I(_0992_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5439_ (.A1(\as2650.stack[3][10] ),
    .A2(_0934_),
    .B(_0937_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5440_ (.I0(\as2650.stack[1][10] ),
    .I1(\as2650.stack[0][10] ),
    .S(_0929_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5441_ (.A1(\as2650.stack[2][10] ),
    .A2(_0920_),
    .B1(_0927_),
    .B2(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5442_ (.A1(_0943_),
    .A2(\as2650.stack[5][10] ),
    .B1(\as2650.stack[4][10] ),
    .B2(_0946_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5443_ (.A1(_0940_),
    .A2(_0997_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5444_ (.A1(_0951_),
    .A2(\as2650.stack[7][10] ),
    .B1(\as2650.stack[6][10] ),
    .B2(_0967_),
    .C(_0973_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5445_ (.A1(_0994_),
    .A2(_0996_),
    .B1(_0998_),
    .B2(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5446_ (.A1(_0993_),
    .A2(_0966_),
    .B1(_1000_),
    .B2(_0982_),
    .C(_0983_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5447_ (.A1(_0396_),
    .A2(_0990_),
    .B(_0991_),
    .C(_1001_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5448_ (.A1(_0988_),
    .A2(_1002_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5449_ (.I(_1003_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5450_ (.A1(\as2650.r123[0][3] ),
    .A2(_0963_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5451_ (.I(_0410_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5452_ (.I(_0921_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5453_ (.I(_1006_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5454_ (.I(_0941_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5455_ (.I(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5456_ (.A1(_1009_),
    .A2(\as2650.stack[5][11] ),
    .B1(\as2650.stack[4][11] ),
    .B2(_0946_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5457_ (.A1(_1007_),
    .A2(_1010_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5458_ (.I(_0950_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5459_ (.A1(_1012_),
    .A2(\as2650.stack[7][11] ),
    .B1(\as2650.stack[6][11] ),
    .B2(_1007_),
    .C(_0954_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5460_ (.I(_0928_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5461_ (.I(_0916_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5462_ (.I0(\as2650.stack[3][11] ),
    .I1(\as2650.stack[0][11] ),
    .I2(\as2650.stack[1][11] ),
    .I3(\as2650.stack[2][11] ),
    .S0(_1014_),
    .S1(_1015_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5463_ (.A1(_0977_),
    .A2(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5464_ (.A1(_1011_),
    .A2(_1013_),
    .B(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5465_ (.I(_0913_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5466_ (.A1(_1005_),
    .A2(_0914_),
    .B1(_1018_),
    .B2(_1019_),
    .C(_0958_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5467_ (.A1(_0987_),
    .A2(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5468_ (.A1(_0493_),
    .A2(_0989_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5469_ (.A1(_1021_),
    .A2(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5470_ (.A1(_1004_),
    .A2(_1023_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5471_ (.A1(\as2650.r123[0][4] ),
    .A2(_0987_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5472_ (.I(_0557_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5473_ (.A1(_0943_),
    .A2(\as2650.stack[5][12] ),
    .B1(\as2650.stack[4][12] ),
    .B2(_0968_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5474_ (.A1(_0967_),
    .A2(_1026_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5475_ (.A1(_0951_),
    .A2(\as2650.stack[7][12] ),
    .B1(\as2650.stack[6][12] ),
    .B2(_0920_),
    .C(_0973_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5476_ (.I0(\as2650.stack[3][12] ),
    .I1(\as2650.stack[0][12] ),
    .I2(\as2650.stack[1][12] ),
    .I3(\as2650.stack[2][12] ),
    .S0(_0929_),
    .S1(_0978_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5477_ (.A1(_0977_),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5478_ (.A1(_1027_),
    .A2(_1028_),
    .B(_1030_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5479_ (.A1(_1025_),
    .A2(_0966_),
    .B1(_1031_),
    .B2(_0982_),
    .C(_0983_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5480_ (.A1(_0599_),
    .A2(_0990_),
    .B(_0991_),
    .C(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5481_ (.A1(_1024_),
    .A2(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5482_ (.I(_1034_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5483_ (.A1(\as2650.r123[0][5] ),
    .A2(_0987_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5484_ (.I(_0655_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5485_ (.I(_0944_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5486_ (.A1(_1009_),
    .A2(\as2650.stack[5][13] ),
    .B1(\as2650.stack[4][13] ),
    .B2(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5487_ (.A1(_0919_),
    .A2(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5488_ (.A1(_1012_),
    .A2(\as2650.stack[7][13] ),
    .B1(\as2650.stack[6][13] ),
    .B2(_1007_),
    .C(_0954_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5489_ (.I0(\as2650.stack[3][13] ),
    .I1(\as2650.stack[0][13] ),
    .I2(\as2650.stack[1][13] ),
    .I3(\as2650.stack[2][13] ),
    .S0(_1014_),
    .S1(_1015_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5490_ (.A1(_0976_),
    .A2(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5491_ (.A1(_1039_),
    .A2(_1040_),
    .B(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5492_ (.A1(_1036_),
    .A2(_0966_),
    .B1(_1043_),
    .B2(_1019_),
    .C(_0983_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5493_ (.A1(_0687_),
    .A2(_0990_),
    .B(_0991_),
    .C(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5494_ (.A1(_1035_),
    .A2(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5495_ (.I(_1046_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5496_ (.A1(\as2650.r123[0][6] ),
    .A2(_0962_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5497_ (.I(_0741_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5498_ (.A1(_1009_),
    .A2(\as2650.stack[5][14] ),
    .B1(\as2650.stack[4][14] ),
    .B2(_0946_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5499_ (.A1(_1007_),
    .A2(_1049_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5500_ (.A1(_1012_),
    .A2(\as2650.stack[7][14] ),
    .B1(\as2650.stack[6][14] ),
    .B2(_0940_),
    .C(_0954_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5501_ (.I0(\as2650.stack[3][14] ),
    .I1(\as2650.stack[0][14] ),
    .I2(\as2650.stack[1][14] ),
    .I3(\as2650.stack[2][14] ),
    .S0(_1014_),
    .S1(_1015_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5502_ (.A1(_0977_),
    .A2(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5503_ (.A1(_1050_),
    .A2(_1051_),
    .B(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5504_ (.A1(_1048_),
    .A2(_0914_),
    .B1(_1054_),
    .B2(_1019_),
    .C(_0958_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5505_ (.A1(_0771_),
    .A2(_0990_),
    .B(_0991_),
    .C(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5506_ (.A1(_1047_),
    .A2(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5507_ (.I(_1057_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5508_ (.A1(\as2650.r123[0][7] ),
    .A2(_0963_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5509_ (.I(_0870_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5510_ (.A1(_1059_),
    .A2(_0957_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5511_ (.A1(_4197_),
    .A2(_0904_),
    .B(_1060_),
    .C(_0894_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5512_ (.A1(_0890_),
    .A2(_0908_),
    .B(_0909_),
    .C(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5513_ (.A1(_1058_),
    .A2(_1062_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5514_ (.I(_0932_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5515_ (.A1(_0335_),
    .A2(_0895_),
    .A3(_0899_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5516_ (.A1(_3934_),
    .A2(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5517_ (.A1(_3905_),
    .A2(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5518_ (.I(_1066_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5519_ (.A1(_0926_),
    .A2(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5520_ (.I(\as2650.halted ),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5521_ (.A1(_1069_),
    .A2(net10),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5522_ (.I(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5523_ (.I(_4007_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5524_ (.I(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5525_ (.A1(_4174_),
    .A2(_0575_),
    .A3(_0911_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5526_ (.A1(_1073_),
    .A2(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5527_ (.A1(_1071_),
    .A2(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5528_ (.A1(_1015_),
    .A2(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5529_ (.A1(_1068_),
    .A2(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5530_ (.A1(_1063_),
    .A2(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5531_ (.A1(_0945_),
    .A2(_1066_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5532_ (.I(_1071_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5533_ (.I(_4204_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5534_ (.A1(_4200_),
    .A2(_4000_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5535_ (.A1(\as2650.ins_reg[3] ),
    .A2(_3958_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5536_ (.A1(_4175_),
    .A2(_1083_),
    .A3(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5537_ (.A1(_1082_),
    .A2(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5538_ (.I(_1086_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5539_ (.I(_3929_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5540_ (.A1(_1088_),
    .A2(_3986_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5541_ (.I(_1089_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5542_ (.I(_1090_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5543_ (.A1(_4154_),
    .A2(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5544_ (.I(\as2650.addr_buff[7] ),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5545_ (.I(_3987_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5546_ (.I(_1094_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5547_ (.I(_3912_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5548_ (.A1(\as2650.cycle[2] ),
    .A2(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5549_ (.A1(\as2650.cycle[3] ),
    .A2(_1088_),
    .A3(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5550_ (.A1(_3955_),
    .A2(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5551_ (.A1(_1093_),
    .A2(_1095_),
    .B(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5552_ (.I(_4170_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5553_ (.I(_3959_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5554_ (.I(_3963_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5555_ (.A1(_4005_),
    .A2(_3943_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5556_ (.A1(_4155_),
    .A2(_4100_),
    .A3(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5557_ (.A1(_1103_),
    .A2(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5558_ (.I(_1106_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5559_ (.A1(_3998_),
    .A2(_1101_),
    .B(_1102_),
    .C(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5560_ (.A1(_4205_),
    .A2(_1100_),
    .B(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5561_ (.A1(_1087_),
    .A2(_1092_),
    .B(_1065_),
    .C(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5562_ (.A1(_1081_),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5563_ (.A1(_1080_),
    .A2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5564_ (.A1(_1079_),
    .A2(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5565_ (.I(_1113_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5566_ (.I(_1114_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5567_ (.I(\as2650.pc[0] ),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5568_ (.I(_1116_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5569_ (.I(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5570_ (.I(_1118_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5571_ (.I0(_4064_),
    .I1(_1119_),
    .S(_1076_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5572_ (.I(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5573_ (.I(_1113_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5574_ (.I(_1122_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5575_ (.A1(\as2650.stack[5][0] ),
    .A2(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5576_ (.A1(_1115_),
    .A2(_1121_),
    .B(_1124_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5577_ (.I(_1067_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5578_ (.I(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5579_ (.I(_1126_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5580_ (.I(\as2650.pc[1] ),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5581_ (.I(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5582_ (.I(_1129_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5583_ (.I(_1125_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5584_ (.A1(_1130_),
    .A2(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5585_ (.A1(_0965_),
    .A2(_1127_),
    .B(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5586_ (.I(_1133_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5587_ (.I(_1122_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5588_ (.A1(\as2650.stack[5][1] ),
    .A2(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5589_ (.A1(_1115_),
    .A2(_1134_),
    .B(_1136_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5590_ (.I(\as2650.pc[2] ),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5591_ (.I(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5592_ (.I(_1138_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5593_ (.A1(_1139_),
    .A2(_1131_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5594_ (.A1(_0993_),
    .A2(_1127_),
    .B(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5595_ (.I(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5596_ (.A1(\as2650.stack[5][2] ),
    .A2(_1135_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5597_ (.A1(_1115_),
    .A2(_1142_),
    .B(_1143_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5598_ (.I(\as2650.pc[3] ),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5599_ (.I(_1144_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5600_ (.A1(_1145_),
    .A2(_1131_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5601_ (.A1(_1005_),
    .A2(_1127_),
    .B(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5602_ (.I(_1147_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5603_ (.A1(\as2650.stack[5][3] ),
    .A2(_1135_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5604_ (.A1(_1115_),
    .A2(_1148_),
    .B(_1149_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5605_ (.I(_1114_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5606_ (.I(\as2650.pc[4] ),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5607_ (.I(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5608_ (.A1(_1152_),
    .A2(_1131_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5609_ (.A1(_1025_),
    .A2(_1127_),
    .B(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5610_ (.I(_1154_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5611_ (.A1(\as2650.stack[5][4] ),
    .A2(_1135_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5612_ (.A1(_1150_),
    .A2(_1155_),
    .B(_1156_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5613_ (.I(_1036_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5614_ (.I(_1126_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5615_ (.I(\as2650.pc[5] ),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5616_ (.I(_1159_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5617_ (.I(_1125_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5618_ (.A1(_1160_),
    .A2(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5619_ (.A1(_1157_),
    .A2(_1158_),
    .B(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5620_ (.I(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5621_ (.I(_1122_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5622_ (.A1(\as2650.stack[5][5] ),
    .A2(_1165_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5623_ (.A1(_1150_),
    .A2(_1164_),
    .B(_1166_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5624_ (.I(_1048_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5625_ (.I(\as2650.pc[6] ),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5626_ (.I(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5627_ (.I(_1169_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5628_ (.A1(_1170_),
    .A2(_1161_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5629_ (.A1(_1167_),
    .A2(_1158_),
    .B(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5630_ (.I(_1172_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5631_ (.A1(\as2650.stack[5][6] ),
    .A2(_1165_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5632_ (.A1(_1150_),
    .A2(_1173_),
    .B(_1174_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5633_ (.I(_0870_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5634_ (.I(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5635_ (.I(\as2650.pc[7] ),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5636_ (.I0(_1176_),
    .I1(_1177_),
    .S(_1076_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5637_ (.I(_1178_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5638_ (.A1(\as2650.stack[5][7] ),
    .A2(_1165_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5639_ (.A1(_1150_),
    .A2(_1179_),
    .B(_1180_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5640_ (.A1(_0953_),
    .A2(_1067_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5641_ (.A1(_1063_),
    .A2(_1067_),
    .B(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5642_ (.A1(_1078_),
    .A2(_1182_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5643_ (.A1(_1081_),
    .A2(_1080_),
    .A3(_1110_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5644_ (.A1(_1183_),
    .A2(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5645_ (.I(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5646_ (.I(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5647_ (.I(\as2650.pc[8] ),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5648_ (.I(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5649_ (.I(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5650_ (.A1(_4223_),
    .A2(_1126_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5651_ (.A1(_1190_),
    .A2(_1076_),
    .B(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5652_ (.I(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5653_ (.I(_1186_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5654_ (.A1(\as2650.stack[6][8] ),
    .A2(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5655_ (.A1(_1187_),
    .A2(_1193_),
    .B(_1195_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5656_ (.I(\as2650.pc[9] ),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5657_ (.I(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5658_ (.I(_1197_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5659_ (.A1(_1198_),
    .A2(_1161_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5660_ (.A1(_0308_),
    .A2(_1158_),
    .B(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5661_ (.I(_1200_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5662_ (.I(_1186_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5663_ (.A1(\as2650.stack[6][9] ),
    .A2(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5664_ (.A1(_1187_),
    .A2(_1201_),
    .B(_1203_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5665_ (.I(\as2650.pc[10] ),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5666_ (.I(_1204_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5667_ (.A1(_1205_),
    .A2(_1161_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5668_ (.A1(_0501_),
    .A2(_1158_),
    .B(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5669_ (.I(_1207_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5670_ (.A1(\as2650.stack[6][10] ),
    .A2(_1202_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5671_ (.A1(_1187_),
    .A2(_1208_),
    .B(_1209_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5672_ (.I(_0831_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5673_ (.I(_1126_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5674_ (.I(\as2650.pc[11] ),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5675_ (.I(_1212_),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5676_ (.I(_1125_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5677_ (.A1(_1213_),
    .A2(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5678_ (.A1(_1210_),
    .A2(_1211_),
    .B(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5679_ (.I(_1216_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5680_ (.A1(\as2650.stack[6][11] ),
    .A2(_1202_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5681_ (.A1(_1187_),
    .A2(_1217_),
    .B(_1218_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5682_ (.I(\as2650.pc[12] ),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5683_ (.I(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5684_ (.I(_1220_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5685_ (.A1(_1221_),
    .A2(_1214_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5686_ (.A1(_0615_),
    .A2(_1211_),
    .B(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5687_ (.I(_1223_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5688_ (.A1(\as2650.stack[6][12] ),
    .A2(_1202_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5689_ (.A1(_1194_),
    .A2(_1224_),
    .B(_1225_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5690_ (.I(\as2650.pc[13] ),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5691_ (.I(_1226_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5692_ (.A1(_1227_),
    .A2(_1214_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5693_ (.A1(_0574_),
    .A2(_1211_),
    .B(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5694_ (.I(_1229_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5695_ (.I(_1186_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5696_ (.A1(\as2650.stack[6][13] ),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5697_ (.A1(_1194_),
    .A2(_1230_),
    .B(_1232_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5698_ (.I(_0786_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5699_ (.I(\as2650.pc[14] ),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5700_ (.A1(_1234_),
    .A2(_1214_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5701_ (.A1(_1233_),
    .A2(_1211_),
    .B(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5702_ (.I(_1236_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5703_ (.A1(\as2650.stack[6][14] ),
    .A2(_1231_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5704_ (.A1(_1194_),
    .A2(_1237_),
    .B(_1238_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5705_ (.I(_3995_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5706_ (.I(_3971_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5707_ (.I(_1093_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5708_ (.A1(_1240_),
    .A2(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5709_ (.I(_3943_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5710_ (.A1(_1096_),
    .A2(_3955_),
    .A3(_3909_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5711_ (.A1(\as2650.cycle[7] ),
    .A2(\as2650.cycle[6] ),
    .A3(_3928_),
    .A4(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5712_ (.A1(_1243_),
    .A2(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5713_ (.I(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5714_ (.A1(_1239_),
    .A2(_4118_),
    .A3(_1242_),
    .B(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5715_ (.I(_1084_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5716_ (.A1(_4025_),
    .A2(_4120_),
    .A3(_4192_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5717_ (.A1(_3900_),
    .A2(_4145_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5718_ (.A1(_1082_),
    .A2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5719_ (.I(_1252_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5720_ (.I(_1103_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5721_ (.I(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5722_ (.I(_1243_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5723_ (.I(_1256_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5724_ (.A1(_1255_),
    .A2(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5725_ (.A1(_1250_),
    .A2(_1253_),
    .A3(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5726_ (.I(_3901_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5727_ (.A1(_1260_),
    .A2(_1073_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5728_ (.A1(_1254_),
    .A2(_1252_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5729_ (.I(_3963_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5730_ (.A1(_1263_),
    .A2(_3961_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5731_ (.A1(_1261_),
    .A2(_1262_),
    .A3(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5732_ (.A1(_1249_),
    .A2(_1259_),
    .A3(_1265_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5733_ (.I(_1094_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5734_ (.I(_1267_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5735_ (.I(_1268_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5736_ (.I(_1072_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_1270_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5738_ (.I(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5739_ (.I(_3960_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5740_ (.A1(_4170_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5741_ (.A1(_1263_),
    .A2(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5742_ (.I(_1275_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5743_ (.A1(_1272_),
    .A2(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5744_ (.I(_1239_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5745_ (.A1(_3951_),
    .A2(_1269_),
    .B1(_1277_),
    .B2(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5746_ (.I(_1069_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5747_ (.I(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5748_ (.A1(_3927_),
    .A2(_3983_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5749_ (.A1(_3982_),
    .A2(_1282_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5750_ (.I(_1283_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5751_ (.I(\as2650.cycle[3] ),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5752_ (.I(_3982_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5753_ (.A1(_1285_),
    .A2(_1286_),
    .A3(_1097_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5754_ (.I(_1287_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5755_ (.A1(_4122_),
    .A2(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5756_ (.A1(_1281_),
    .A2(_4186_),
    .A3(_1284_),
    .A4(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5757_ (.I(_3934_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5758_ (.A1(_1260_),
    .A2(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5759_ (.I(_1292_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5760_ (.I(_1282_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5761_ (.A1(_3911_),
    .A2(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5762_ (.A1(_3907_),
    .A2(_1295_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5763_ (.I(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5764_ (.A1(_4121_),
    .A2(_1283_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5765_ (.I(net3),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5766_ (.I(_1299_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5767_ (.I(_1300_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5768_ (.I(\as2650.cycle[6] ),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5769_ (.A1(\as2650.cycle[7] ),
    .A2(_3910_),
    .A3(_1282_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5770_ (.A1(_1302_),
    .A2(_1303_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5771_ (.A1(_1301_),
    .A2(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5772_ (.A1(_1293_),
    .A2(_1297_),
    .B1(_1298_),
    .B2(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5773_ (.A1(_1290_),
    .A2(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5774_ (.A1(_1248_),
    .A2(_1266_),
    .A3(_1279_),
    .A4(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5775_ (.A1(_3909_),
    .A2(_3982_),
    .A3(_3973_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5776_ (.I(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5777_ (.I(_1245_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5778_ (.A1(_1311_),
    .A2(_1090_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5779_ (.A1(_1292_),
    .A2(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5780_ (.A1(_3971_),
    .A2(_3910_),
    .A3(_1294_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5781_ (.A1(_1302_),
    .A2(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5782_ (.A1(_1313_),
    .A2(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5783_ (.A1(_1310_),
    .A2(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5784_ (.A1(_1243_),
    .A2(_4008_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5785_ (.A1(_3956_),
    .A2(_3987_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5786_ (.A1(_1318_),
    .A2(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5787_ (.A1(_3907_),
    .A2(_3915_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5788_ (.A1(_1321_),
    .A2(_1296_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5789_ (.A1(_1287_),
    .A2(_1303_),
    .A3(_1320_),
    .A4(_1322_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5790_ (.A1(_3975_),
    .A2(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5791_ (.A1(_1308_),
    .A2(_1317_),
    .A3(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5792_ (.I(_1325_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5793_ (.I(_1239_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5794_ (.A1(_1327_),
    .A2(_3920_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5795_ (.I(_1328_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5796_ (.I(_1328_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5797_ (.A1(_4064_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5798_ (.A1(_0872_),
    .A2(_1329_),
    .B(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5799_ (.I(_1325_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5800_ (.A1(net41),
    .A2(_1333_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5801_ (.A1(_1326_),
    .A2(_1332_),
    .B(_1334_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5802_ (.I(_0350_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5803_ (.A1(_1335_),
    .A2(_1330_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5804_ (.A1(_0965_),
    .A2(_1329_),
    .B(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5805_ (.A1(net42),
    .A2(_1333_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5806_ (.A1(_1326_),
    .A2(_1337_),
    .B(_1338_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5807_ (.I(_1328_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5808_ (.I(_1328_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5809_ (.A1(_0442_),
    .A2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5810_ (.A1(_0993_),
    .A2(_1339_),
    .B(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5811_ (.A1(net43),
    .A2(_1333_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5812_ (.A1(_1326_),
    .A2(_1342_),
    .B(_1343_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5813_ (.I(_0410_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5814_ (.I(_0523_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5815_ (.A1(_1345_),
    .A2(_1340_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5816_ (.A1(_1344_),
    .A2(_1339_),
    .B(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5817_ (.A1(net44),
    .A2(_1333_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5818_ (.A1(_1326_),
    .A2(_1347_),
    .B(_1348_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5819_ (.I(_1325_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5820_ (.I(_0557_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5821_ (.I(_0422_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5822_ (.A1(_1351_),
    .A2(_1340_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5823_ (.A1(_1350_),
    .A2(_1339_),
    .B(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5824_ (.I(_1325_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5825_ (.A1(net45),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5826_ (.A1(_1349_),
    .A2(_1353_),
    .B(_1355_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5827_ (.I(_0639_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5828_ (.A1(_1356_),
    .A2(_1340_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5829_ (.A1(_1157_),
    .A2(_1339_),
    .B(_1357_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5830_ (.A1(net19),
    .A2(_1354_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5831_ (.A1(_1349_),
    .A2(_1358_),
    .B(_1359_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5832_ (.I(_0676_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5833_ (.I(_1360_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5834_ (.I(_0741_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5835_ (.A1(_1362_),
    .A2(_1330_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5836_ (.A1(_1361_),
    .A2(_1329_),
    .B(_1363_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5837_ (.A1(net20),
    .A2(_1354_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5838_ (.A1(_1349_),
    .A2(_1364_),
    .B(_1365_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5839_ (.A1(_1176_),
    .A2(_1330_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5840_ (.A1(_4107_),
    .A2(_1329_),
    .B(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5841_ (.A1(net21),
    .A2(_1354_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5842_ (.A1(_1349_),
    .A2(_1367_),
    .B(_1368_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5843_ (.I(\as2650.psu[5] ),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5844_ (.I(_1253_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5845_ (.I(_4025_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5846_ (.A1(_1371_),
    .A2(_0660_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5847_ (.A1(_1372_),
    .A2(_4029_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5848_ (.A1(_1273_),
    .A2(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5849_ (.I(_1374_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5850_ (.I(_4009_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5851_ (.A1(_4196_),
    .A2(_0901_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5852_ (.A1(_4200_),
    .A2(_0892_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5853_ (.A1(_4174_),
    .A2(_4195_),
    .A3(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5854_ (.I(_3991_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5855_ (.A1(_0906_),
    .A2(_1380_),
    .A3(_0911_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5856_ (.A1(_1074_),
    .A2(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5857_ (.A1(_1376_),
    .A2(_1377_),
    .A3(_1379_),
    .A4(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5858_ (.A1(_1370_),
    .A2(_1375_),
    .A3(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5859_ (.I(_0438_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5860_ (.A1(_3991_),
    .A2(_1378_),
    .A3(_0910_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5861_ (.I(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5862_ (.I(_1387_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5863_ (.I(_0902_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5864_ (.A1(_4196_),
    .A2(_1389_),
    .A3(_1074_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5865_ (.I(_1083_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5866_ (.A1(_4009_),
    .A2(_0851_),
    .A3(_1391_),
    .A4(_0899_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5867_ (.A1(_1385_),
    .A2(_1388_),
    .B(_1390_),
    .C(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5868_ (.A1(_3934_),
    .A2(_1245_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5869_ (.I(_1394_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5870_ (.I(_1395_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5871_ (.I(_4100_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5872_ (.A1(\as2650.psl[6] ),
    .A2(_3999_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5873_ (.A1(\as2650.psl[7] ),
    .A2(_4000_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5874_ (.A1(_1398_),
    .A2(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5875_ (.A1(_1397_),
    .A2(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5876_ (.A1(_1271_),
    .A2(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5877_ (.A1(_0538_),
    .A2(_1402_),
    .B(_1370_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5878_ (.A1(_4204_),
    .A2(_4005_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5879_ (.A1(_1102_),
    .A2(_4027_),
    .A3(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5880_ (.I(_1405_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5881_ (.A1(_1253_),
    .A2(_1375_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5882_ (.I(_3956_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5883_ (.I(_1408_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5884_ (.I(_1409_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5885_ (.A1(_1391_),
    .A2(_1406_),
    .B(_1407_),
    .C(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5886_ (.I(_4006_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5887_ (.I(_1412_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5888_ (.I(_1413_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5889_ (.I(_1245_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5890_ (.I(_4204_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5891_ (.A1(_1416_),
    .A2(_4006_),
    .A3(_3997_),
    .A4(_4203_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5892_ (.A1(_0895_),
    .A2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5893_ (.A1(_1415_),
    .A2(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5894_ (.A1(_1280_),
    .A2(_1309_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5895_ (.I(_1420_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5896_ (.A1(_1414_),
    .A2(_1375_),
    .A3(_1419_),
    .A4(_1421_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5897_ (.A1(_1396_),
    .A2(_1403_),
    .A3(_1411_),
    .A4(_1422_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5898_ (.A1(_1384_),
    .A2(_1393_),
    .A3(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5899_ (.I(_1370_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5900_ (.A1(_1036_),
    .A2(_1385_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5901_ (.I(_0658_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5902_ (.I(_1427_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5903_ (.I(_1270_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5904_ (.I(_1429_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5905_ (.I(_1430_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5906_ (.A1(_4003_),
    .A2(_1417_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5907_ (.A1(_1427_),
    .A2(_1432_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5908_ (.A1(\as2650.psu[5] ),
    .A2(_1428_),
    .B(_1431_),
    .C(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5909_ (.A1(_1426_),
    .A2(_1434_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5910_ (.A1(_1425_),
    .A2(_1435_),
    .B(_1424_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5911_ (.I(_4187_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5912_ (.I(_1437_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5913_ (.A1(_1369_),
    .A2(_1424_),
    .B(_1436_),
    .C(_1438_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5914_ (.I(\as2650.r123_2[3][0] ),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5915_ (.I(_1439_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5916_ (.I(\as2650.r123_2[3][1] ),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5917_ (.I(_1440_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5918_ (.I(\as2650.r123_2[3][2] ),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5919_ (.I(_1441_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5920_ (.I(\as2650.r123_2[3][3] ),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5921_ (.I(_1442_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5922_ (.I(\as2650.r123_2[3][4] ),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5923_ (.I(_1443_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5924_ (.I(\as2650.r123_2[3][5] ),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5925_ (.I(_1444_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5926_ (.I(\as2650.r123_2[3][6] ),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5927_ (.I(_1445_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5928_ (.I(\as2650.r123_2[3][7] ),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5929_ (.I(_1446_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5930_ (.A1(_1012_),
    .A2(_1078_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5931_ (.A1(_1184_),
    .A2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5932_ (.I(_1448_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5933_ (.I(_1449_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5934_ (.I(_1448_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5935_ (.I(_1451_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5936_ (.A1(\as2650.stack[0][8] ),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5937_ (.A1(_1193_),
    .A2(_1450_),
    .B(_1453_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5938_ (.I(_1451_),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5939_ (.A1(\as2650.stack[0][9] ),
    .A2(_1454_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5940_ (.A1(_1201_),
    .A2(_1450_),
    .B(_1455_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5941_ (.A1(\as2650.stack[0][10] ),
    .A2(_1454_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5942_ (.A1(_1208_),
    .A2(_1450_),
    .B(_1456_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5943_ (.A1(\as2650.stack[0][11] ),
    .A2(_1454_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5944_ (.A1(_1217_),
    .A2(_1450_),
    .B(_1457_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5945_ (.I(_1449_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5946_ (.A1(\as2650.stack[0][12] ),
    .A2(_1454_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5947_ (.A1(_1224_),
    .A2(_1458_),
    .B(_1459_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5948_ (.I(_1451_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5949_ (.A1(\as2650.stack[0][13] ),
    .A2(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5950_ (.A1(_1230_),
    .A2(_1458_),
    .B(_1461_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5951_ (.A1(\as2650.stack[0][14] ),
    .A2(_1460_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5952_ (.A1(_1237_),
    .A2(_1458_),
    .B(_1462_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5953_ (.A1(_1112_),
    .A2(_1447_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5954_ (.I(_1463_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5955_ (.I(_1464_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5956_ (.I(_1463_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5957_ (.I(_1466_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5958_ (.A1(\as2650.stack[1][8] ),
    .A2(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5959_ (.A1(_1193_),
    .A2(_1465_),
    .B(_1468_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5960_ (.I(_1466_),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5961_ (.A1(\as2650.stack[1][9] ),
    .A2(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5962_ (.A1(_1201_),
    .A2(_1465_),
    .B(_1470_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5963_ (.A1(\as2650.stack[1][10] ),
    .A2(_1469_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5964_ (.A1(_1208_),
    .A2(_1465_),
    .B(_1471_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5965_ (.A1(\as2650.stack[1][11] ),
    .A2(_1469_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5966_ (.A1(_1217_),
    .A2(_1465_),
    .B(_1472_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5967_ (.I(_1464_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5968_ (.A1(\as2650.stack[1][12] ),
    .A2(_1469_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5969_ (.A1(_1224_),
    .A2(_1473_),
    .B(_1474_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5970_ (.I(_1466_),
    .Z(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5971_ (.A1(\as2650.stack[1][13] ),
    .A2(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5972_ (.A1(_1230_),
    .A2(_1473_),
    .B(_1476_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5973_ (.A1(\as2650.stack[1][14] ),
    .A2(_1475_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5974_ (.A1(_1237_),
    .A2(_1473_),
    .B(_1477_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5975_ (.I(_1192_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5976_ (.A1(_1068_),
    .A2(_1077_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5977_ (.A1(_1479_),
    .A2(_1182_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5978_ (.A1(_1184_),
    .A2(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5979_ (.I(_1481_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5980_ (.I(_1482_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5981_ (.I(_1481_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5982_ (.I(_1484_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5983_ (.A1(\as2650.stack[2][8] ),
    .A2(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5984_ (.A1(_1478_),
    .A2(_1483_),
    .B(_1486_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5985_ (.I(_1200_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5986_ (.I(_1484_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5987_ (.A1(\as2650.stack[2][9] ),
    .A2(_1488_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5988_ (.A1(_1487_),
    .A2(_1483_),
    .B(_1489_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5989_ (.I(_1207_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5990_ (.A1(\as2650.stack[2][10] ),
    .A2(_1488_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5991_ (.A1(_1490_),
    .A2(_1483_),
    .B(_1491_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5992_ (.I(_1216_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5993_ (.A1(\as2650.stack[2][11] ),
    .A2(_1488_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5994_ (.A1(_1492_),
    .A2(_1483_),
    .B(_1493_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5995_ (.I(_1223_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5996_ (.I(_1482_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5997_ (.A1(\as2650.stack[2][12] ),
    .A2(_1488_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5998_ (.A1(_1494_),
    .A2(_1495_),
    .B(_1496_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5999_ (.I(_1229_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6000_ (.I(_1484_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6001_ (.A1(\as2650.stack[2][13] ),
    .A2(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6002_ (.A1(_1497_),
    .A2(_1495_),
    .B(_1499_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6003_ (.I(_1236_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6004_ (.A1(\as2650.stack[2][14] ),
    .A2(_1498_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6005_ (.A1(_1500_),
    .A2(_1495_),
    .B(_1501_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6006_ (.I(_0845_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6007_ (.I(_4174_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6008_ (.A1(_0856_),
    .A2(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6009_ (.A1(_1503_),
    .A2(_0738_),
    .B(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6010_ (.A1(_0522_),
    .A2(_0630_),
    .A3(_0845_),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6011_ (.A1(_0532_),
    .A2(_0754_),
    .A3(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6012_ (.A1(_0857_),
    .A2(_1505_),
    .B(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6013_ (.A1(\as2650.psl[1] ),
    .A2(_1502_),
    .B(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6014_ (.A1(_0519_),
    .A2(_0539_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6015_ (.A1(_1510_),
    .A2(_0760_),
    .B(_0761_),
    .C(_0751_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6016_ (.A1(_0750_),
    .A2(_1502_),
    .A3(_1511_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6017_ (.A1(\as2650.psl[1] ),
    .A2(_1502_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6018_ (.I(_1505_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6019_ (.A1(_1513_),
    .A2(_1514_),
    .B(_4280_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6020_ (.A1(_1509_),
    .A2(_1512_),
    .A3(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6021_ (.I(_1516_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6022_ (.I(_0769_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6023_ (.A1(_4183_),
    .A2(_0301_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6024_ (.A1(_0348_),
    .A2(_0491_),
    .A3(_0547_),
    .A4(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6025_ (.A1(_0647_),
    .A2(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6026_ (.A1(_4280_),
    .A2(_0861_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6027_ (.A1(_1518_),
    .A2(_1521_),
    .B(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6028_ (.I(_1293_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6029_ (.I(_1524_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6030_ (.A1(_1517_),
    .A2(_1523_),
    .B(_1525_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6031_ (.I(_3961_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6032_ (.I(_1527_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6033_ (.I(_1528_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6034_ (.I(_4070_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6035_ (.I(_4272_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6036_ (.I(_0353_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6037_ (.I(_0427_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6038_ (.A1(_1530_),
    .A2(_1531_),
    .A3(_1532_),
    .A4(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6039_ (.I(_0561_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6040_ (.I(net2),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6041_ (.I(_1536_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6042_ (.I(_1537_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6043_ (.I(_1538_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6044_ (.I(_1539_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6045_ (.I(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6046_ (.A1(_1535_),
    .A2(_1427_),
    .A3(_1541_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6047_ (.I(_0876_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6048_ (.I(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6049_ (.A1(_1534_),
    .A2(_1542_),
    .B(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6050_ (.A1(_1416_),
    .A2(_1256_),
    .A3(_4292_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6051_ (.A1(_1546_),
    .A2(_0873_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6052_ (.I(_0738_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6053_ (.A1(_1335_),
    .A2(_1548_),
    .A3(_0445_),
    .A4(_0865_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6054_ (.I(_1527_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6055_ (.A1(_0374_),
    .A2(_4246_),
    .A3(_4214_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6056_ (.A1(_0741_),
    .A2(_0655_),
    .A3(_0417_),
    .A4(_0366_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6057_ (.A1(_1551_),
    .A2(_1552_),
    .B(_0869_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6058_ (.A1(_1362_),
    .A2(_1381_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6059_ (.I(_1291_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6060_ (.I(_1555_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6061_ (.A1(_1381_),
    .A2(_1553_),
    .B(_1554_),
    .C(_1556_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6062_ (.A1(\as2650.psl[6] ),
    .A2(_1539_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6063_ (.A1(_0892_),
    .A2(_1540_),
    .B(_1558_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6064_ (.A1(_4202_),
    .A2(_1430_),
    .A3(_1406_),
    .A4(_1559_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6065_ (.I(_4020_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6066_ (.A1(_1557_),
    .A2(_1560_),
    .B(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6067_ (.I(_1372_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6068_ (.I(_1563_),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6069_ (.A1(_4110_),
    .A2(_0718_),
    .B(_1361_),
    .C(_1564_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6070_ (.I(_4029_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6071_ (.I(_1566_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6072_ (.A1(_1562_),
    .A2(_1565_),
    .B(_1567_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6073_ (.A1(_1547_),
    .A2(_1549_),
    .B(_1550_),
    .C(_1568_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6074_ (.I(_1278_),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6075_ (.I(_1570_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6076_ (.A1(_1529_),
    .A2(_1545_),
    .B(_1569_),
    .C(_1571_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6077_ (.I(_1410_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6078_ (.A1(_1391_),
    .A2(_1406_),
    .B(_1407_),
    .C(_1573_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6079_ (.I(_4005_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6080_ (.A1(_1575_),
    .A2(_1260_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6081_ (.I(_1576_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6082_ (.A1(_0538_),
    .A2(_1577_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6083_ (.A1(_1103_),
    .A2(_0436_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6084_ (.A1(_1546_),
    .A2(_1579_),
    .B(_1275_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6085_ (.I(_1408_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6086_ (.A1(_4201_),
    .A2(_1581_),
    .A3(_1417_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6087_ (.A1(_1320_),
    .A2(_1390_),
    .A3(_1582_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6088_ (.A1(_1580_),
    .A2(_1583_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6089_ (.A1(_1380_),
    .A2(_4195_),
    .A3(_0575_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6090_ (.A1(_4145_),
    .A2(_1576_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6091_ (.A1(_4196_),
    .A2(_1585_),
    .A3(_1375_),
    .A4(_1586_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6092_ (.A1(_3991_),
    .A2(_4195_),
    .A3(_1397_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6093_ (.A1(_1383_),
    .A2(_1588_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6094_ (.A1(_1587_),
    .A2(_1589_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6095_ (.I(_1311_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6096_ (.A1(_3957_),
    .A2(_1251_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6097_ (.I(_1592_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6098_ (.A1(_1263_),
    .A2(_1593_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6099_ (.A1(_4122_),
    .A2(_1376_),
    .A3(_1594_),
    .A4(_1374_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6100_ (.A1(_1591_),
    .A2(_1595_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6101_ (.A1(_4024_),
    .A2(_3952_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6102_ (.I(_1597_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6103_ (.I(_4015_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6104_ (.A1(_0851_),
    .A2(_1261_),
    .B1(_1598_),
    .B2(_1599_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6105_ (.A1(_4020_),
    .A2(_1579_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6106_ (.A1(_1264_),
    .A2(_1395_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6107_ (.A1(_1600_),
    .A2(_1601_),
    .A3(_1602_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6108_ (.A1(_1380_),
    .A2(_4203_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6109_ (.A1(_1243_),
    .A2(_4191_),
    .A3(_4148_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6110_ (.A1(_1072_),
    .A2(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6111_ (.A1(_1069_),
    .A2(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6112_ (.A1(_1247_),
    .A2(_1607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6113_ (.A1(_0436_),
    .A2(_1379_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6114_ (.A1(_1104_),
    .A2(_1593_),
    .A3(_1608_),
    .A4(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6115_ (.A1(_1088_),
    .A2(_1294_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6116_ (.A1(_3972_),
    .A2(_1088_),
    .A3(_3973_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6117_ (.A1(_1611_),
    .A2(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6118_ (.A1(_1260_),
    .A2(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6119_ (.A1(_1257_),
    .A2(_0898_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6120_ (.A1(_4015_),
    .A2(_1605_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6121_ (.A1(_0850_),
    .A2(_1598_),
    .A3(_1616_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6122_ (.A1(_3952_),
    .A2(_1614_),
    .A3(_1615_),
    .A4(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6123_ (.A1(_1272_),
    .A2(_1604_),
    .B(_1610_),
    .C(_1618_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6124_ (.A1(_1590_),
    .A2(_1596_),
    .A3(_1603_),
    .A4(_1619_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6125_ (.A1(_1574_),
    .A2(_1578_),
    .B(_1584_),
    .C(_1620_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6126_ (.I(_1261_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6127_ (.I(_1622_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6128_ (.I(_1548_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6129_ (.A1(_1257_),
    .A2(_0898_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6130_ (.I(_1625_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6131_ (.A1(_1624_),
    .A2(_0866_),
    .A3(_1626_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6132_ (.A1(_1553_),
    .A2(_1615_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6133_ (.A1(_1627_),
    .A2(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6134_ (.A1(_1623_),
    .A2(_1629_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6135_ (.A1(_1526_),
    .A2(_1572_),
    .A3(_1621_),
    .A4(_1630_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6136_ (.I(_3903_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6137_ (.I(_1632_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6138_ (.A1(\as2650.psl[6] ),
    .A2(_1621_),
    .B(_1633_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6139_ (.A1(_1631_),
    .A2(_1634_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6140_ (.I(_1632_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6141_ (.I(\as2650.psl[7] ),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6142_ (.A1(_4289_),
    .A2(_0296_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6143_ (.A1(_0754_),
    .A2(_1506_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6144_ (.A1(_4142_),
    .A2(_0529_),
    .A3(_1637_),
    .A4(_1638_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6145_ (.A1(_4280_),
    .A2(_1639_),
    .B(_1522_),
    .C(_1516_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6146_ (.A1(_1548_),
    .A2(_1626_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6147_ (.A1(_1059_),
    .A2(_1626_),
    .B(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6148_ (.A1(_1101_),
    .A2(_1250_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6149_ (.A1(_1527_),
    .A2(_1547_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6150_ (.I(_1599_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6151_ (.A1(_0869_),
    .A2(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6152_ (.I(_0874_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6153_ (.A1(_1397_),
    .A2(_1405_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6154_ (.A1(_4175_),
    .A2(_1102_),
    .A3(_1404_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6155_ (.A1(_3885_),
    .A2(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6156_ (.I(\as2650.psu[3] ),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6157_ (.I(net1),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6158_ (.A1(_0935_),
    .A2(_4270_),
    .B1(_0352_),
    .B2(_0932_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6159_ (.A1(\as2650.psu[7] ),
    .A2(_1299_),
    .B1(_1652_),
    .B2(\as2650.psu[5] ),
    .C(_1653_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6160_ (.I(_0558_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6161_ (.I(_4069_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _6162_ (.A1(\as2650.psu[4] ),
    .A2(_1655_),
    .B1(_0729_),
    .B2(net27),
    .C1(_0915_),
    .C2(_1656_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6163_ (.A1(_1651_),
    .A2(_0425_),
    .B(_1654_),
    .C(_1657_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6164_ (.A1(_1650_),
    .A2(_1658_),
    .B(_1648_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6165_ (.I(_1655_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6166_ (.I(\as2650.psl[3] ),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6167_ (.I(_0351_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6168_ (.I(_1662_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6169_ (.A1(\as2650.psl[7] ),
    .A2(_1299_),
    .B1(_1663_),
    .B2(\as2650.overflow ),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6170_ (.A1(_4108_),
    .A2(_4069_),
    .B1(_0424_),
    .B2(_1661_),
    .C(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6171_ (.I(\as2650.psl[1] ),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6172_ (.I(\as2650.psl[5] ),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6173_ (.I(\as2650.psl[6] ),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6174_ (.A1(_1666_),
    .A2(_4270_),
    .B1(_0656_),
    .B2(_1667_),
    .C1(_1537_),
    .C2(_1668_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6175_ (.A1(_3969_),
    .A2(_1660_),
    .B(_1665_),
    .C(_1669_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6176_ (.A1(_4201_),
    .A2(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6177_ (.A1(_0874_),
    .A2(_0737_),
    .B1(_0442_),
    .B2(_0352_),
    .C1(_0639_),
    .C2(_0657_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6178_ (.I(_1656_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6179_ (.I(_0559_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6180_ (.A1(_4269_),
    .A2(_0295_),
    .B1(_0421_),
    .B2(_1674_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6181_ (.A1(_1673_),
    .A2(_0871_),
    .B1(_0675_),
    .B2(_0729_),
    .C(_1675_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6182_ (.A1(_0425_),
    .A2(_0523_),
    .B1(_1649_),
    .B2(_4201_),
    .C(_1676_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6183_ (.A1(_1649_),
    .A2(_1671_),
    .B1(_1672_),
    .B2(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6184_ (.A1(_1636_),
    .A2(_1647_),
    .A3(_1648_),
    .B1(_1659_),
    .B2(_1678_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6185_ (.A1(_1418_),
    .A2(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6186_ (.A1(_1636_),
    .A2(_1301_),
    .A3(_1418_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6187_ (.A1(_1680_),
    .A2(_1681_),
    .B(_1429_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6188_ (.A1(_1646_),
    .A2(_1682_),
    .B(_0439_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6189_ (.I(_1546_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6190_ (.A1(_1561_),
    .A2(_1360_),
    .B(_1683_),
    .C(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6191_ (.A1(_1644_),
    .A2(_1685_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6192_ (.I(_1256_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6193_ (.I(_1687_),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6194_ (.A1(_1544_),
    .A2(_1643_),
    .B(_1686_),
    .C(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6195_ (.A1(_1524_),
    .A2(_1640_),
    .B1(_1642_),
    .B2(_1622_),
    .C(_1689_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6196_ (.I0(_1636_),
    .I1(_1690_),
    .S(_1621_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6197_ (.A1(_1635_),
    .A2(_1691_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6198_ (.I(_1692_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6199_ (.A1(\as2650.stack[0][0] ),
    .A2(_1460_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6200_ (.A1(_1121_),
    .A2(_1458_),
    .B(_1693_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6201_ (.I(_1451_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6202_ (.A1(\as2650.stack[0][1] ),
    .A2(_1460_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6203_ (.A1(_1134_),
    .A2(_1694_),
    .B(_1695_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6204_ (.I(_1448_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6205_ (.A1(\as2650.stack[0][2] ),
    .A2(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6206_ (.A1(_1142_),
    .A2(_1694_),
    .B(_1697_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6207_ (.A1(\as2650.stack[0][3] ),
    .A2(_1696_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6208_ (.A1(_1148_),
    .A2(_1694_),
    .B(_1698_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6209_ (.A1(\as2650.stack[0][4] ),
    .A2(_1696_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6210_ (.A1(_1155_),
    .A2(_1694_),
    .B(_1699_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6211_ (.A1(\as2650.stack[0][5] ),
    .A2(_1696_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6212_ (.A1(_1164_),
    .A2(_1452_),
    .B(_1700_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6213_ (.A1(\as2650.stack[0][6] ),
    .A2(_1449_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6214_ (.A1(_1173_),
    .A2(_1452_),
    .B(_1701_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6215_ (.A1(\as2650.stack[0][7] ),
    .A2(_1449_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6216_ (.A1(_1179_),
    .A2(_1452_),
    .B(_1702_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6217_ (.A1(\as2650.stack[1][0] ),
    .A2(_1475_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6218_ (.A1(_1121_),
    .A2(_1473_),
    .B(_1703_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6219_ (.I(_1466_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6220_ (.A1(\as2650.stack[1][1] ),
    .A2(_1475_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6221_ (.A1(_1134_),
    .A2(_1704_),
    .B(_1705_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6222_ (.I(_1463_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6223_ (.A1(\as2650.stack[1][2] ),
    .A2(_1706_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6224_ (.A1(_1142_),
    .A2(_1704_),
    .B(_1707_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6225_ (.A1(\as2650.stack[1][3] ),
    .A2(_1706_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6226_ (.A1(_1148_),
    .A2(_1704_),
    .B(_1708_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6227_ (.A1(\as2650.stack[1][4] ),
    .A2(_1706_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6228_ (.A1(_1155_),
    .A2(_1704_),
    .B(_1709_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6229_ (.A1(\as2650.stack[1][5] ),
    .A2(_1706_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6230_ (.A1(_1164_),
    .A2(_1467_),
    .B(_1710_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6231_ (.A1(\as2650.stack[1][6] ),
    .A2(_1464_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6232_ (.A1(_1173_),
    .A2(_1467_),
    .B(_1711_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(\as2650.stack[1][7] ),
    .A2(_1464_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6234_ (.A1(_1179_),
    .A2(_1467_),
    .B(_1712_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6235_ (.A1(_1371_),
    .A2(_1085_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6236_ (.A1(_1300_),
    .A2(_1408_),
    .A3(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6237_ (.A1(_1310_),
    .A2(_1714_),
    .B(_1081_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6238_ (.I(_1715_),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6239_ (.I(_1530_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6240_ (.I(_1310_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6241_ (.I(_1715_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6242_ (.I(_1249_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6243_ (.I(_1720_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6244_ (.A1(_1721_),
    .A2(_1310_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6245_ (.A1(_1717_),
    .A2(_1718_),
    .B(_1719_),
    .C(_1722_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6246_ (.A1(_3885_),
    .A2(_1716_),
    .B(_1723_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6247_ (.A1(_1531_),
    .A2(_1718_),
    .B(_1719_),
    .C(_1722_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6248_ (.A1(_0892_),
    .A2(_1716_),
    .B(_1724_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6249_ (.I(_0353_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6250_ (.A1(_4037_),
    .A2(_1612_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6251_ (.I(_1726_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6252_ (.I(_1416_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6253_ (.I(_1728_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6254_ (.A1(_1725_),
    .A2(_1727_),
    .B1(_1716_),
    .B2(_1729_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6255_ (.I(_1730_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6256_ (.I(_1105_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6257_ (.A1(_1416_),
    .A2(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6258_ (.I(_1732_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6259_ (.I(_1733_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6260_ (.I(_1734_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6261_ (.I(_1735_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6262_ (.A1(_4164_),
    .A2(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6263_ (.A1(_1428_),
    .A2(_1718_),
    .B1(_1722_),
    .B2(_1737_),
    .C(_1715_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6264_ (.A1(_4164_),
    .A2(_1716_),
    .B(_1738_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6265_ (.I(_1541_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6266_ (.A1(_1739_),
    .A2(_1727_),
    .B1(_1719_),
    .B2(_3998_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6267_ (.I(_1740_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6268_ (.I(_1543_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6269_ (.A1(_1741_),
    .A2(_1726_),
    .B1(_1719_),
    .B2(_1101_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6270_ (.I(_1742_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6271_ (.A1(\as2650.stack[2][0] ),
    .A2(_1498_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6272_ (.A1(_1121_),
    .A2(_1495_),
    .B(_1743_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6273_ (.I(_1484_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6274_ (.A1(\as2650.stack[2][1] ),
    .A2(_1498_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6275_ (.A1(_1134_),
    .A2(_1744_),
    .B(_1745_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6276_ (.I(_1481_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6277_ (.A1(\as2650.stack[2][2] ),
    .A2(_1746_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6278_ (.A1(_1142_),
    .A2(_1744_),
    .B(_1747_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6279_ (.A1(\as2650.stack[2][3] ),
    .A2(_1746_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6280_ (.A1(_1148_),
    .A2(_1744_),
    .B(_1748_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6281_ (.A1(\as2650.stack[2][4] ),
    .A2(_1746_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6282_ (.A1(_1155_),
    .A2(_1744_),
    .B(_1749_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6283_ (.A1(\as2650.stack[2][5] ),
    .A2(_1746_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6284_ (.A1(_1164_),
    .A2(_1485_),
    .B(_1750_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6285_ (.A1(\as2650.stack[2][6] ),
    .A2(_1482_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6286_ (.A1(_1173_),
    .A2(_1485_),
    .B(_1751_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6287_ (.A1(\as2650.stack[2][7] ),
    .A2(_1482_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6288_ (.A1(_1179_),
    .A2(_1485_),
    .B(_1752_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6289_ (.A1(_1112_),
    .A2(_1480_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6290_ (.I(_1753_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6291_ (.I(_1754_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6292_ (.I(_1753_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6293_ (.I(_1756_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6294_ (.A1(\as2650.stack[3][8] ),
    .A2(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6295_ (.A1(_1478_),
    .A2(_1755_),
    .B(_1758_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6296_ (.I(_1756_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6297_ (.A1(\as2650.stack[3][9] ),
    .A2(_1759_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6298_ (.A1(_1487_),
    .A2(_1755_),
    .B(_1760_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6299_ (.A1(\as2650.stack[3][10] ),
    .A2(_1759_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6300_ (.A1(_1490_),
    .A2(_1755_),
    .B(_1761_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6301_ (.A1(\as2650.stack[3][11] ),
    .A2(_1759_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6302_ (.A1(_1492_),
    .A2(_1755_),
    .B(_1762_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6303_ (.I(_1754_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6304_ (.A1(\as2650.stack[3][12] ),
    .A2(_1759_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6305_ (.A1(_1494_),
    .A2(_1763_),
    .B(_1764_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6306_ (.I(_1756_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6307_ (.A1(\as2650.stack[3][13] ),
    .A2(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6308_ (.A1(_1497_),
    .A2(_1763_),
    .B(_1766_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6309_ (.A1(\as2650.stack[3][14] ),
    .A2(_1765_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6310_ (.A1(_1500_),
    .A2(_1763_),
    .B(_1767_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6311_ (.A1(_3969_),
    .A2(_1071_),
    .A3(_4015_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6312_ (.A1(_4197_),
    .A2(_1768_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6313_ (.I(_1769_),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6314_ (.I(_1770_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6315_ (.A1(_0812_),
    .A2(_0841_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6316_ (.A1(_0809_),
    .A2(_0842_),
    .B(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6317_ (.A1(_0818_),
    .A2(_0839_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6318_ (.A1(_0815_),
    .A2(_0840_),
    .B(_1774_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6319_ (.A1(_0869_),
    .A2(_4222_),
    .A3(_0835_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6320_ (.A1(_0832_),
    .A2(_0837_),
    .B(_1776_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6321_ (.A1(_0823_),
    .A2(_0829_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6322_ (.A1(_0823_),
    .A2(_0829_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6323_ (.A1(_0819_),
    .A2(_1778_),
    .A3(_1779_),
    .B1(_0830_),
    .B2(_0838_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6324_ (.A1(_0666_),
    .A2(_0306_),
    .A3(_0822_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6325_ (.A1(_0796_),
    .A2(_0821_),
    .B(_1781_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6326_ (.A1(_0580_),
    .A2(_0831_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6327_ (.A1(_1782_),
    .A2(_1783_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6328_ (.A1(_0789_),
    .A2(_0828_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6329_ (.A1(_0823_),
    .A2(_0829_),
    .B(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6330_ (.A1(\as2650.r0[7] ),
    .A2(_0304_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6331_ (.A1(\as2650.r0[6] ),
    .A2(\as2650.r0[4] ),
    .A3(_0399_),
    .A4(_0611_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6332_ (.A1(\as2650.r0[6] ),
    .A2(_0400_),
    .B1(_0612_),
    .B2(_0414_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6333_ (.A1(_1788_),
    .A2(_1789_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6334_ (.A1(_1787_),
    .A2(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6335_ (.I(_0826_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6336_ (.A1(_0497_),
    .A2(_1792_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6337_ (.A1(_0824_),
    .A2(_0827_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6338_ (.A1(_0787_),
    .A2(_1793_),
    .B1(_1794_),
    .B2(_0825_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6339_ (.A1(_0364_),
    .A2(_0788_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6340_ (.A1(_4254_),
    .A2(_0786_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6341_ (.A1(_1793_),
    .A2(_1796_),
    .A3(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6342_ (.A1(_1791_),
    .A2(_1795_),
    .A3(_1798_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6343_ (.A1(_1786_),
    .A2(_1799_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6344_ (.A1(_1784_),
    .A2(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6345_ (.A1(_1780_),
    .A2(_1801_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6346_ (.A1(_1777_),
    .A2(_1802_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6347_ (.A1(_1773_),
    .A2(_1775_),
    .A3(_1803_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6348_ (.A1(_1771_),
    .A2(_1804_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6349_ (.I(_3936_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6350_ (.A1(_1806_),
    .A2(_3952_),
    .A3(_1768_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6351_ (.I(_1807_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6352_ (.A1(_3925_),
    .A2(_1070_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6353_ (.A1(_4008_),
    .A2(_1809_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6354_ (.A1(_4024_),
    .A2(_4030_),
    .A3(_1810_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6355_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6356_ (.A1(_3925_),
    .A2(_4002_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6357_ (.A1(_4040_),
    .A2(_1813_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6358_ (.I(_1814_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6359_ (.I(_1809_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6360_ (.A1(_3993_),
    .A2(_1816_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6361_ (.A1(_3890_),
    .A2(_4001_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6362_ (.I(_1818_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6363_ (.A1(_3962_),
    .A2(_3965_),
    .A3(_1819_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6364_ (.I(_1820_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6365_ (.A1(_4014_),
    .A2(_3964_),
    .A3(_4019_),
    .A4(_1818_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6366_ (.I(_1822_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6367_ (.A1(_3975_),
    .A2(_3979_),
    .A3(_1813_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6368_ (.A1(_1821_),
    .A2(_1823_),
    .A3(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6369_ (.A1(_4011_),
    .A2(_1816_),
    .B(_1817_),
    .C(_1825_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6370_ (.A1(_1808_),
    .A2(_1812_),
    .A3(_1815_),
    .A4(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6371_ (.A1(_1391_),
    .A2(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6372_ (.A1(_1770_),
    .A2(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6373_ (.I(_1829_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6374_ (.A1(_0495_),
    .A2(_1810_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6375_ (.A1(_3994_),
    .A2(_1816_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6376_ (.I(_1832_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6377_ (.A1(_3923_),
    .A2(_1819_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6378_ (.I(_1834_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6379_ (.A1(_4119_),
    .A2(_4124_),
    .A3(_1819_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6380_ (.I(_1836_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6381_ (.A1(_4003_),
    .A2(_1503_),
    .A3(_3951_),
    .A4(_1810_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6382_ (.I(_1838_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6383_ (.A1(_4214_),
    .A2(_1839_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6384_ (.I(_4095_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6385_ (.A1(_1841_),
    .A2(_1548_),
    .B(_4161_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6386_ (.I(_1822_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6387_ (.I(_1843_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6388_ (.I(_1823_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6389_ (.A1(_4206_),
    .A2(_1813_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6390_ (.I(_1846_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6391_ (.A1(_1412_),
    .A2(_1071_),
    .A3(_3962_),
    .A4(_1819_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6392_ (.A1(_0659_),
    .A2(_4251_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6393_ (.I(_1811_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6394_ (.A1(_4070_),
    .A2(_1847_),
    .B1(_1848_),
    .B2(_1849_),
    .C(_1850_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6395_ (.A1(_0350_),
    .A2(_1812_),
    .B(_1845_),
    .C(_1851_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6396_ (.I(_1807_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6397_ (.A1(_1842_),
    .A2(_1844_),
    .B(_1852_),
    .C(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6398_ (.A1(_1840_),
    .A2(_1854_),
    .B(_1835_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6399_ (.A1(_4062_),
    .A2(_1835_),
    .B(_1837_),
    .C(_1855_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6400_ (.I(_1824_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6401_ (.I(_1857_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6402_ (.A1(_4131_),
    .A2(_1858_),
    .B(_1832_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6403_ (.A1(_4183_),
    .A2(_1833_),
    .B1(_1856_),
    .B2(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6404_ (.A1(_1831_),
    .A2(_1860_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6405_ (.I(_1828_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6406_ (.A1(\as2650.r123_2[2][0] ),
    .A2(_1830_),
    .B1(_1861_),
    .B2(_1862_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6407_ (.A1(_1805_),
    .A2(_1863_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6408_ (.A1(_1775_),
    .A2(_1803_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6409_ (.A1(_1775_),
    .A2(_1803_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6410_ (.A1(_1773_),
    .A2(_1864_),
    .B(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6411_ (.A1(_1780_),
    .A2(_1801_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6412_ (.A1(_1777_),
    .A2(_1802_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6413_ (.A1(_1867_),
    .A2(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6414_ (.A1(_0655_),
    .A2(_1210_),
    .A3(_1782_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6415_ (.A1(_1786_),
    .A2(_1799_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6416_ (.A1(_1784_),
    .A2(_1800_),
    .B(_1871_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6417_ (.A1(_1787_),
    .A2(_1790_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6418_ (.A1(_1788_),
    .A2(_1873_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6419_ (.A1(_0665_),
    .A2(_0505_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6420_ (.A1(_1874_),
    .A2(_1875_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6421_ (.A1(_1795_),
    .A2(_1798_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6422_ (.A1(_1795_),
    .A2(_1798_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6423_ (.A1(_1791_),
    .A2(_1877_),
    .B(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6424_ (.A1(_4096_),
    .A2(_0403_),
    .B1(_0614_),
    .B2(_0580_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6425_ (.A1(_4096_),
    .A2(_0614_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6426_ (.A1(_0821_),
    .A2(_1881_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6427_ (.A1(_1880_),
    .A2(_1882_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6428_ (.A1(_4254_),
    .A2(_0826_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6429_ (.A1(_1793_),
    .A2(_1797_),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6430_ (.A1(_0824_),
    .A2(_1884_),
    .B1(_1885_),
    .B2(_1796_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6431_ (.A1(_0415_),
    .A2(_0788_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6432_ (.A1(\as2650.r0[3] ),
    .A2(_0785_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6433_ (.A1(_1884_),
    .A2(_1888_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6434_ (.A1(_1887_),
    .A2(_1889_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6435_ (.A1(_1886_),
    .A2(_1890_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6436_ (.A1(_1883_),
    .A2(_1891_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6437_ (.A1(_1876_),
    .A2(_1879_),
    .A3(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6438_ (.A1(_1872_),
    .A2(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6439_ (.A1(_1870_),
    .A2(_1894_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6440_ (.A1(_1869_),
    .A2(_1895_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6441_ (.A1(_1866_),
    .A2(_1896_),
    .Z(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6442_ (.A1(_1771_),
    .A2(_1897_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6443_ (.I(_1769_),
    .Z(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6444_ (.I(_1814_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6445_ (.A1(_4271_),
    .A2(_1821_),
    .B(_1850_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6446_ (.A1(_4267_),
    .A2(_1847_),
    .B(_1901_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6447_ (.I(_1811_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6448_ (.A1(_0442_),
    .A2(_1903_),
    .B(_1843_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6449_ (.A1(_0872_),
    .A2(_1844_),
    .B1(_1902_),
    .B2(_1904_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6450_ (.A1(_1853_),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6451_ (.A1(_4246_),
    .A2(_1853_),
    .B(_1900_),
    .C(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6452_ (.A1(_4244_),
    .A2(_1835_),
    .B(_1837_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6453_ (.A1(_4236_),
    .A2(_1837_),
    .B1(_1907_),
    .B2(_1908_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6454_ (.I(_1832_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6455_ (.A1(_0301_),
    .A2(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6456_ (.A1(_1833_),
    .A2(_1909_),
    .B(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6457_ (.A1(_1899_),
    .A2(_1912_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6458_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_1830_),
    .B1(_1913_),
    .B2(_1862_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6459_ (.A1(_1898_),
    .A2(_1914_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6460_ (.A1(_1869_),
    .A2(_1895_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6461_ (.A1(_1866_),
    .A2(_1896_),
    .B(_1915_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6462_ (.A1(_1872_),
    .A2(_1893_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6463_ (.A1(_1870_),
    .A2(_1894_),
    .B(_1917_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6464_ (.A1(_1874_),
    .A2(_1875_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6465_ (.A1(_1879_),
    .A2(_1892_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6466_ (.A1(_1879_),
    .A2(_1892_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6467_ (.A1(_1876_),
    .A2(_1920_),
    .B(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6468_ (.A1(_1210_),
    .A2(_1882_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6469_ (.A1(_4096_),
    .A2(_0831_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6470_ (.A1(_0821_),
    .A2(_1881_),
    .B(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6471_ (.A1(_1923_),
    .A2(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6472_ (.A1(_1886_),
    .A2(_1890_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6473_ (.A1(_1883_),
    .A2(_1891_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6474_ (.A1(_1927_),
    .A2(_1928_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6475_ (.A1(_0665_),
    .A2(_0614_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6476_ (.A1(\as2650.r0[3] ),
    .A2(_0826_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6477_ (.A1(_1797_),
    .A2(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6478_ (.A1(_1887_),
    .A2(_1889_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6479_ (.A1(_1932_),
    .A2(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6480_ (.A1(\as2650.r0[4] ),
    .A2(_0784_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6481_ (.A1(_1931_),
    .A2(_1935_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6482_ (.A1(_0579_),
    .A2(_0788_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6483_ (.A1(_1936_),
    .A2(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6484_ (.A1(_1934_),
    .A2(_1938_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6485_ (.A1(_1930_),
    .A2(_1939_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6486_ (.A1(_1929_),
    .A2(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6487_ (.A1(_1926_),
    .A2(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6488_ (.A1(_1922_),
    .A2(_1942_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6489_ (.A1(_1919_),
    .A2(_1943_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6490_ (.A1(_1918_),
    .A2(_1944_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6491_ (.A1(_1916_),
    .A2(_1945_),
    .Z(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6492_ (.A1(_1771_),
    .A2(_1946_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6493_ (.I(_1829_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6494_ (.I(_1769_),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6495_ (.I(_1817_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6496_ (.I(_1824_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6497_ (.I(_1823_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6498_ (.A1(_4260_),
    .A2(_0358_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6499_ (.I(_1662_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6500_ (.A1(_1954_),
    .A2(_1820_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6501_ (.A1(_4003_),
    .A2(_4030_),
    .A3(_1810_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6502_ (.A1(_1953_),
    .A2(_1846_),
    .B(_1955_),
    .C(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6503_ (.A1(_0370_),
    .A2(_1850_),
    .B(_1823_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6504_ (.A1(_0350_),
    .A2(_1952_),
    .B1(_1957_),
    .B2(_1958_),
    .C(_1807_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6505_ (.A1(_0374_),
    .A2(_1808_),
    .B(_1815_),
    .C(_1959_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6506_ (.A1(_0386_),
    .A2(_1815_),
    .B(_1857_),
    .C(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6507_ (.A1(_0393_),
    .A2(_1951_),
    .B(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6508_ (.A1(_1950_),
    .A2(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6509_ (.A1(_0349_),
    .A2(_1950_),
    .B(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6510_ (.A1(_1949_),
    .A2(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6511_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_1948_),
    .B1(_1965_),
    .B2(_1862_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6512_ (.A1(_1947_),
    .A2(_1966_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6513_ (.A1(_1918_),
    .A2(_1944_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6514_ (.A1(_1916_),
    .A2(_1945_),
    .B(_1967_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6515_ (.I(_1943_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6516_ (.A1(_1922_),
    .A2(_1942_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6517_ (.A1(_1919_),
    .A2(_1969_),
    .B(_1970_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6518_ (.A1(_0416_),
    .A2(_1792_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6519_ (.A1(_1888_),
    .A2(_1972_),
    .B1(_1936_),
    .B2(_1937_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6520_ (.A1(_0579_),
    .A2(_0786_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6521_ (.A1(_1972_),
    .A2(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6522_ (.A1(_0666_),
    .A2(_0573_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6523_ (.A1(_1975_),
    .A2(_1976_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6524_ (.A1(_1973_),
    .A2(_1977_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6525_ (.A1(_1881_),
    .A2(_1978_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6526_ (.A1(_0667_),
    .A2(_0615_),
    .A3(_1939_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6527_ (.A1(_1934_),
    .A2(_1938_),
    .B(_1980_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6528_ (.A1(_1979_),
    .A2(_1981_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6529_ (.I(_1940_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6530_ (.A1(_1929_),
    .A2(_1983_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6531_ (.A1(_1923_),
    .A2(_1925_),
    .A3(_1941_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6532_ (.A1(_1984_),
    .A2(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6533_ (.A1(_1982_),
    .A2(_1986_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6534_ (.A1(_1923_),
    .A2(_1987_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6535_ (.A1(_1968_),
    .A2(_1971_),
    .A3(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6536_ (.A1(_1771_),
    .A2(_1989_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6537_ (.A1(_0426_),
    .A2(_1821_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6538_ (.A1(_0433_),
    .A2(_1821_),
    .B(_1991_),
    .C(_1956_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6539_ (.A1(_0422_),
    .A2(_1903_),
    .B(_1843_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6540_ (.A1(_4260_),
    .A2(_1845_),
    .B1(_1992_),
    .B2(_1993_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6541_ (.I(_1838_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6542_ (.A1(_0410_),
    .A2(_1995_),
    .B(_1834_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6543_ (.A1(_1839_),
    .A2(_1994_),
    .B(_1996_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6544_ (.A1(_0454_),
    .A2(_1900_),
    .B(_1857_),
    .C(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6545_ (.A1(_0460_),
    .A2(_1858_),
    .B(_1998_),
    .C(_1832_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6546_ (.A1(_0492_),
    .A2(_1833_),
    .B(_1999_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6547_ (.A1(_1899_),
    .A2(_2000_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6548_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_1948_),
    .B1(_2001_),
    .B2(_1862_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6549_ (.A1(_1990_),
    .A2(_2002_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6550_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_1830_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6551_ (.A1(_1982_),
    .A2(_1986_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6552_ (.A1(_1923_),
    .A2(_1987_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6553_ (.A1(_1979_),
    .A2(_1981_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6554_ (.A1(_0580_),
    .A2(_1792_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6555_ (.A1(_1935_),
    .A2(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6556_ (.A1(_1975_),
    .A2(_1976_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6557_ (.A1(_2008_),
    .A2(_2009_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6558_ (.A1(_0666_),
    .A2(_1233_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6559_ (.A1(_2007_),
    .A2(_2011_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6560_ (.A1(_4097_),
    .A2(_0574_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6561_ (.A1(_2012_),
    .A2(_2013_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6562_ (.A1(_2010_),
    .A2(_2014_),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6563_ (.A1(_2010_),
    .A2(_2014_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6564_ (.A1(_2015_),
    .A2(_2016_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6565_ (.I(_1973_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6566_ (.A1(_1881_),
    .A2(_1978_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6567_ (.A1(_2018_),
    .A2(_1977_),
    .B(_2019_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6568_ (.A1(_2017_),
    .A2(_2020_),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6569_ (.A1(_2006_),
    .A2(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6570_ (.A1(_2004_),
    .A2(_2005_),
    .B(_2022_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6571_ (.A1(_2004_),
    .A2(_2005_),
    .A3(_2022_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6572_ (.A1(_2023_),
    .A2(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6573_ (.A1(_1971_),
    .A2(_1988_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6574_ (.A1(_1971_),
    .A2(_1988_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6575_ (.A1(_1968_),
    .A2(_2026_),
    .B(_2027_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6576_ (.A1(_2025_),
    .A2(_2028_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6577_ (.A1(_0557_),
    .A2(_1995_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6578_ (.I(_0560_),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6579_ (.A1(_0564_),
    .A2(_1846_),
    .B(_1956_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6580_ (.A1(_2031_),
    .A2(_1846_),
    .B(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6581_ (.A1(_1356_),
    .A2(_1903_),
    .B(_1952_),
    .C(_2033_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6582_ (.A1(_0370_),
    .A2(_1844_),
    .B(_2034_),
    .C(_1808_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6583_ (.I(_1834_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6584_ (.A1(_2030_),
    .A2(_2035_),
    .B(_2036_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6585_ (.A1(_0594_),
    .A2(_1835_),
    .B(_1837_),
    .C(_2037_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6586_ (.A1(_0556_),
    .A2(_1951_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6587_ (.A1(_1950_),
    .A2(_2038_),
    .A3(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6588_ (.A1(_0548_),
    .A2(_1950_),
    .B(_2040_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6589_ (.A1(_1899_),
    .A2(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6590_ (.I(_1828_),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6591_ (.A1(_1949_),
    .A2(_2029_),
    .B1(_2042_),
    .B2(_2043_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6592_ (.A1(_2003_),
    .A2(_2044_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6593_ (.A1(_2025_),
    .A2(_2028_),
    .B(_2023_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6594_ (.A1(_2006_),
    .A2(_2021_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6595_ (.I(_2017_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6596_ (.A1(_2047_),
    .A2(_2020_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6597_ (.A1(_2015_),
    .A2(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6598_ (.I(_1792_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6599_ (.A1(_0667_),
    .A2(_2050_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6600_ (.A1(_1974_),
    .A2(_2051_),
    .B1(_2012_),
    .B2(_2013_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6601_ (.A1(_4097_),
    .A2(_1233_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6602_ (.A1(_2051_),
    .A2(_2053_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6603_ (.A1(_2052_),
    .A2(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6604_ (.A1(_2049_),
    .A2(_2055_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6605_ (.A1(_2046_),
    .A2(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6606_ (.A1(_2045_),
    .A2(_2057_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6607_ (.A1(_1949_),
    .A2(_2058_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6608_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_1830_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6609_ (.I(_1831_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6610_ (.I(_0648_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6611_ (.I(_1652_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6612_ (.A1(_2063_),
    .A2(_1847_),
    .B1(_1848_),
    .B2(_0662_),
    .C(_1850_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6613_ (.A1(_1360_),
    .A2(_1812_),
    .B(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6614_ (.A1(_0544_),
    .A2(_1845_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6615_ (.A1(_1844_),
    .A2(_2065_),
    .B(_2066_),
    .C(_1995_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6616_ (.A1(_1036_),
    .A2(_1839_),
    .B(_2036_),
    .C(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6617_ (.A1(_0682_),
    .A2(_1900_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6618_ (.A1(_2068_),
    .A2(_2069_),
    .B(_1951_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6619_ (.A1(_0654_),
    .A2(_1858_),
    .B(_2070_),
    .C(_1910_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6620_ (.A1(_2062_),
    .A2(_1833_),
    .B(_2071_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6621_ (.A1(_2061_),
    .A2(_2043_),
    .A3(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6622_ (.A1(_2059_),
    .A2(_2060_),
    .A3(_2073_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6623_ (.I(_2061_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6624_ (.A1(_2046_),
    .A2(_2056_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6625_ (.A1(_2045_),
    .A2(_2057_),
    .B(_2075_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6626_ (.A1(_2048_),
    .A2(_2055_),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6627_ (.A1(_0870_),
    .A2(_2050_),
    .A3(_2011_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6628_ (.A1(_2052_),
    .A2(_2054_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6629_ (.A1(_2015_),
    .A2(_2055_),
    .B(_2079_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6630_ (.A1(_2078_),
    .A2(_2080_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6631_ (.A1(_2076_),
    .A2(_2077_),
    .A3(_2081_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6632_ (.I(_0728_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6633_ (.I(_2083_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6634_ (.A1(_2084_),
    .A2(_1820_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6635_ (.A1(_1956_),
    .A2(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6636_ (.A1(_0733_),
    .A2(_1848_),
    .B(_2086_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6637_ (.A1(_0738_),
    .A2(_1812_),
    .B(_1952_),
    .C(_2087_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6638_ (.A1(_0586_),
    .A2(_1952_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6639_ (.A1(_1995_),
    .A2(_2089_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6640_ (.A1(_1048_),
    .A2(_1839_),
    .B1(_2088_),
    .B2(_2090_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6641_ (.A1(_0726_),
    .A2(_2036_),
    .B(_1836_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6642_ (.A1(_2036_),
    .A2(_2091_),
    .B(_2092_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6643_ (.A1(_0722_),
    .A2(_1951_),
    .B(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6644_ (.I0(_0769_),
    .I1(_2094_),
    .S(_1817_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6645_ (.A1(_1899_),
    .A2(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6646_ (.A1(\as2650.r123_2[2][6] ),
    .A2(_1948_),
    .B1(_2096_),
    .B2(_2043_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6647_ (.A1(_2074_),
    .A2(_2082_),
    .B(_2097_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6648_ (.A1(_2077_),
    .A2(_2081_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6649_ (.I(_2080_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6650_ (.A1(_1059_),
    .A2(_2050_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6651_ (.A1(_2011_),
    .A2(_2099_),
    .B(_2100_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6652_ (.A1(_2077_),
    .A2(_2081_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6653_ (.A1(_2076_),
    .A2(_2098_),
    .B(_2101_),
    .C(_2102_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6654_ (.I(_0868_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6655_ (.A1(_1647_),
    .A2(_1820_),
    .B(_1811_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6656_ (.A1(_0878_),
    .A2(_1847_),
    .B(_2105_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6657_ (.A1(_0873_),
    .A2(_1903_),
    .B(_1843_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6658_ (.A1(_1360_),
    .A2(_1845_),
    .B1(_2106_),
    .B2(_2107_),
    .C(_1808_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6659_ (.A1(_1175_),
    .A2(_1853_),
    .B(_1815_),
    .C(_2108_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6660_ (.A1(_0886_),
    .A2(_1900_),
    .B(_1857_),
    .C(_2109_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6661_ (.A1(_2104_),
    .A2(_1858_),
    .B(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6662_ (.A1(_0861_),
    .A2(_1910_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6663_ (.A1(_1910_),
    .A2(_2111_),
    .B(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6664_ (.A1(_1770_),
    .A2(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6665_ (.A1(\as2650.r123_2[2][7] ),
    .A2(_1948_),
    .B1(_2114_),
    .B2(_2043_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6666_ (.A1(_2061_),
    .A2(_2103_),
    .B(_2115_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6667_ (.I(_1120_),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6668_ (.A1(_1079_),
    .A2(_1184_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6669_ (.I(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6670_ (.I(_2118_),
    .Z(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6671_ (.I(_2117_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6672_ (.I(_2120_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6673_ (.A1(\as2650.stack[4][0] ),
    .A2(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6674_ (.A1(_2116_),
    .A2(_2119_),
    .B(_2122_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6675_ (.I(_1133_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6676_ (.I(_2120_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6677_ (.A1(\as2650.stack[4][1] ),
    .A2(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6678_ (.A1(_2123_),
    .A2(_2119_),
    .B(_2125_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6679_ (.I(_1141_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6680_ (.A1(\as2650.stack[4][2] ),
    .A2(_2124_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6681_ (.A1(_2126_),
    .A2(_2119_),
    .B(_2127_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6682_ (.I(_1147_),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6683_ (.A1(\as2650.stack[4][3] ),
    .A2(_2124_),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6684_ (.A1(_2128_),
    .A2(_2119_),
    .B(_2129_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6685_ (.I(_1154_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6686_ (.I(_2118_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6687_ (.A1(\as2650.stack[4][4] ),
    .A2(_2124_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6688_ (.A1(_2130_),
    .A2(_2131_),
    .B(_2132_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6689_ (.I(_1163_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6690_ (.I(_2120_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6691_ (.A1(\as2650.stack[4][5] ),
    .A2(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6692_ (.A1(_2133_),
    .A2(_2131_),
    .B(_2135_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6693_ (.I(_1172_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6694_ (.A1(\as2650.stack[4][6] ),
    .A2(_2134_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6695_ (.A1(_2136_),
    .A2(_2131_),
    .B(_2137_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6696_ (.I(_1178_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6697_ (.A1(\as2650.stack[4][7] ),
    .A2(_2134_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6698_ (.A1(_2138_),
    .A2(_2131_),
    .B(_2139_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6699_ (.A1(\as2650.stack[3][0] ),
    .A2(_1765_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6700_ (.A1(_2116_),
    .A2(_1763_),
    .B(_2140_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6701_ (.I(_1756_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6702_ (.A1(\as2650.stack[3][1] ),
    .A2(_1765_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6703_ (.A1(_2123_),
    .A2(_2141_),
    .B(_2142_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6704_ (.I(_1753_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6705_ (.A1(\as2650.stack[3][2] ),
    .A2(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6706_ (.A1(_2126_),
    .A2(_2141_),
    .B(_2144_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6707_ (.A1(\as2650.stack[3][3] ),
    .A2(_2143_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6708_ (.A1(_2128_),
    .A2(_2141_),
    .B(_2145_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6709_ (.A1(\as2650.stack[3][4] ),
    .A2(_2143_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6710_ (.A1(_2130_),
    .A2(_2141_),
    .B(_2146_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6711_ (.A1(\as2650.stack[3][5] ),
    .A2(_2143_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6712_ (.A1(_2133_),
    .A2(_1757_),
    .B(_2147_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6713_ (.A1(\as2650.stack[3][6] ),
    .A2(_1754_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6714_ (.A1(_2136_),
    .A2(_1757_),
    .B(_2148_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6715_ (.A1(\as2650.stack[3][7] ),
    .A2(_1754_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6716_ (.A1(_2138_),
    .A2(_1757_),
    .B(_2149_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6717_ (.A1(_0906_),
    .A2(_1827_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6718_ (.I(_2150_),
    .Z(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6719_ (.A1(_1860_),
    .A2(_2151_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6720_ (.A1(_1389_),
    .A2(_1768_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6721_ (.A1(_2150_),
    .A2(_2153_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6722_ (.A1(\as2650.r123_2[0][0] ),
    .A2(_2154_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6723_ (.I(_0900_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6724_ (.I(_2156_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6725_ (.A1(_1073_),
    .A2(_0912_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6726_ (.I(_2158_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6727_ (.A1(_4036_),
    .A2(_1081_),
    .A3(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6728_ (.I(_2153_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6729_ (.A1(_2157_),
    .A2(_0956_),
    .B1(_2160_),
    .B2(_4216_),
    .C(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6730_ (.A1(_2152_),
    .A2(_2155_),
    .A3(_2162_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6731_ (.A1(_0906_),
    .A2(_1827_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6732_ (.I(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6733_ (.I(_2154_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6734_ (.I(_2153_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6735_ (.A1(_2157_),
    .A2(_0981_),
    .B1(_2160_),
    .B2(_0310_),
    .C(_2166_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6736_ (.I(_2167_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6737_ (.A1(\as2650.r123_2[0][1] ),
    .A2(_2165_),
    .B(_2168_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6738_ (.A1(_1912_),
    .A2(_2164_),
    .B(_2169_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6739_ (.A1(_1555_),
    .A2(_0900_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6740_ (.A1(_2170_),
    .A2(_1816_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6741_ (.A1(_0992_),
    .A2(_1019_),
    .B1(_1000_),
    .B2(_2171_),
    .C(_2166_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6742_ (.I(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6743_ (.A1(\as2650.r123_2[0][2] ),
    .A2(_2165_),
    .B(_2173_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6744_ (.A1(_1964_),
    .A2(_2164_),
    .B(_2174_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6745_ (.A1(_2157_),
    .A2(_1018_),
    .B1(_2160_),
    .B2(_1005_),
    .C(_2166_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6746_ (.I(_2175_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6747_ (.A1(\as2650.r123_2[0][3] ),
    .A2(_2165_),
    .B(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6748_ (.A1(_2000_),
    .A2(_2164_),
    .B(_2177_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6749_ (.A1(_2157_),
    .A2(_1031_),
    .B1(_2160_),
    .B2(_1025_),
    .C(_2166_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6750_ (.I(_2178_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6751_ (.A1(\as2650.r123_2[0][4] ),
    .A2(_2165_),
    .B(_2179_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6752_ (.A1(_2041_),
    .A2(_2164_),
    .B(_2180_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6753_ (.A1(_2072_),
    .A2(_2151_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6754_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_2154_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6755_ (.A1(_1157_),
    .A2(_0982_),
    .B1(_1043_),
    .B2(_2171_),
    .C(_2161_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6756_ (.A1(_2181_),
    .A2(_2182_),
    .A3(_2183_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6757_ (.A1(_1048_),
    .A2(_0957_),
    .B1(_1054_),
    .B2(_2171_),
    .C(_2153_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6758_ (.I(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6759_ (.A1(\as2650.r123_2[0][6] ),
    .A2(_2154_),
    .B(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6760_ (.A1(_2095_),
    .A2(_2163_),
    .B(_2186_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6761_ (.A1(\as2650.r123_2[0][7] ),
    .A2(_2151_),
    .A3(_2161_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6762_ (.A1(_2113_),
    .A2(_2151_),
    .B1(_2161_),
    .B2(_1060_),
    .C(_2187_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6763_ (.I(_1770_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6764_ (.A1(_4216_),
    .A2(_4223_),
    .A3(_2188_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6765_ (.A1(_4202_),
    .A2(_1827_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6766_ (.I(_2190_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6767_ (.A1(_1769_),
    .A2(_2190_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6768_ (.I(_2192_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6769_ (.A1(_1861_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(\as2650.r123_2[1][0] ),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6770_ (.A1(_2189_),
    .A2(_2194_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6771_ (.I(_2192_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6772_ (.A1(_1913_),
    .A2(_2191_),
    .B1(_2195_),
    .B2(\as2650.r123_2[1][1] ),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6773_ (.A1(_0313_),
    .A2(_2074_),
    .B(_2196_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6774_ (.I(_2190_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6775_ (.A1(_1965_),
    .A2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6776_ (.A1(_0407_),
    .A2(_2188_),
    .B1(_2193_),
    .B2(\as2650.r123_2[1][2] ),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6777_ (.A1(_2198_),
    .A2(_2199_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6778_ (.A1(_2001_),
    .A2(_2191_),
    .B1(_2195_),
    .B2(\as2650.r123_2[1][3] ),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6779_ (.A1(_0513_),
    .A2(_2074_),
    .B(_2200_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6780_ (.A1(_2042_),
    .A2(_2197_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6781_ (.A1(_0624_),
    .A2(_2188_),
    .B1(_2193_),
    .B2(\as2650.r123_2[1][4] ),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6782_ (.A1(_2201_),
    .A2(_2202_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6783_ (.A1(_2061_),
    .A2(_2072_),
    .A3(_2197_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6784_ (.A1(_0712_),
    .A2(_2188_),
    .B1(_2193_),
    .B2(\as2650.r123_2[1][5] ),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6785_ (.A1(_2203_),
    .A2(_2204_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6786_ (.A1(_2096_),
    .A2(_2197_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6787_ (.A1(_0806_),
    .A2(_1949_),
    .B1(_2195_),
    .B2(\as2650.r123_2[1][6] ),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6788_ (.A1(_2205_),
    .A2(_2206_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6789_ (.A1(_2114_),
    .A2(_2191_),
    .B1(_2195_),
    .B2(\as2650.r123_2[1][7] ),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6790_ (.A1(_0843_),
    .A2(_2074_),
    .B(_2207_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6791_ (.I(\as2650.r123[3][0] ),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6792_ (.I(_2208_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6793_ (.I(\as2650.r123[3][1] ),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6794_ (.I(_2209_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6795_ (.I(\as2650.r123[3][2] ),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6796_ (.I(_2210_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6797_ (.I(\as2650.r123[3][3] ),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6798_ (.I(_2211_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6799_ (.I(\as2650.r123[3][4] ),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6800_ (.I(_2212_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6801_ (.I(\as2650.r123[3][5] ),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6802_ (.I(_2213_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6803_ (.I(\as2650.r123[3][6] ),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6804_ (.I(_2214_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6805_ (.I(\as2650.r123[3][7] ),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6806_ (.I(_2215_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6807_ (.I(_3917_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6808_ (.I(_1581_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6809_ (.A1(_2216_),
    .A2(_2217_),
    .A3(_1293_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6810_ (.I(_0437_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6811_ (.A1(_1371_),
    .A2(_1731_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6812_ (.A1(_3913_),
    .A2(_1098_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6813_ (.A1(_1094_),
    .A2(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6814_ (.A1(_1311_),
    .A2(_1084_),
    .A3(_2220_),
    .A4(_2222_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6815_ (.A1(_2219_),
    .A2(_1734_),
    .A3(_2223_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6816_ (.A1(_1249_),
    .A2(_2218_),
    .B(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6817_ (.A1(_1073_),
    .A2(_1107_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6818_ (.I(_1095_),
    .Z(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6819_ (.I(_2227_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6820_ (.I(_1713_),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6821_ (.A1(_2228_),
    .A2(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6822_ (.I(_1104_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6823_ (.A1(_1278_),
    .A2(_2226_),
    .B1(_2230_),
    .B2(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6824_ (.A1(_1280_),
    .A2(net10),
    .A3(_1284_),
    .A4(_1289_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6825_ (.A1(_4121_),
    .A2(_1304_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6826_ (.I(_3973_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6827_ (.A1(_1286_),
    .A2(_2235_),
    .A3(_3985_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6828_ (.A1(_1409_),
    .A2(_1267_),
    .A3(_2220_),
    .A4(_2236_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6829_ (.A1(_4279_),
    .A2(_1309_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6830_ (.I(_1731_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6831_ (.A1(_1082_),
    .A2(_1084_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6832_ (.A1(_1376_),
    .A2(_1311_),
    .A3(_2239_),
    .A4(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6833_ (.A1(_2237_),
    .A2(_2238_),
    .A3(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6834_ (.A1(_2233_),
    .A2(_1323_),
    .A3(_2234_),
    .A4(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6835_ (.A1(_2225_),
    .A2(_2232_),
    .A3(_2243_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6836_ (.I(_2244_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6837_ (.I(_2245_),
    .Z(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6838_ (.I(\as2650.addr_buff[0] ),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6839_ (.I(_2244_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6840_ (.A1(_2247_),
    .A2(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6841_ (.A1(_1673_),
    .A2(_2246_),
    .B(_2249_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6842_ (.I(_4268_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6843_ (.I(_2250_),
    .Z(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6844_ (.I(\as2650.addr_buff[1] ),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6845_ (.I(_2244_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6846_ (.A1(_2252_),
    .A2(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6847_ (.A1(_2251_),
    .A2(_2246_),
    .B(_2254_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6848_ (.I(_1954_),
    .Z(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6849_ (.I(\as2650.addr_buff[2] ),
    .Z(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6850_ (.A1(_2256_),
    .A2(_2253_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6851_ (.A1(_2255_),
    .A2(_2246_),
    .B(_2257_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6852_ (.I(_1533_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6853_ (.I(\as2650.addr_buff[3] ),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6854_ (.I0(_2258_),
    .I1(_2259_),
    .S(_2245_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6855_ (.I(_2260_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6856_ (.I(\as2650.addr_buff[4] ),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6857_ (.A1(_2261_),
    .A2(_2253_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6858_ (.A1(_1660_),
    .A2(_2246_),
    .B(_2262_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6859_ (.I(_3919_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6860_ (.A1(_2263_),
    .A2(_2253_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6861_ (.A1(_2063_),
    .A2(_2248_),
    .B(_2264_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6862_ (.I(_3918_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6863_ (.A1(_2265_),
    .A2(_2245_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6864_ (.A1(_0730_),
    .A2(_2248_),
    .B(_2266_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6865_ (.I(_1301_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6866_ (.I(_1241_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6867_ (.A1(_2268_),
    .A2(_2245_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6868_ (.A1(_2267_),
    .A2(_2248_),
    .B(_2269_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6869_ (.A1(_1413_),
    .A2(_1253_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6870_ (.I(_2270_),
    .Z(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6871_ (.I(_1274_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6872_ (.I(_1645_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6873_ (.A1(_3949_),
    .A2(_1250_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6874_ (.A1(_2273_),
    .A2(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6875_ (.A1(_1247_),
    .A2(_1421_),
    .A3(_2238_),
    .A4(_2275_),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6876_ (.A1(_2271_),
    .A2(_2272_),
    .A3(_1319_),
    .B(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6877_ (.A1(_1288_),
    .A2(_1320_),
    .B(_2277_),
    .C(_1266_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6878_ (.I(_1327_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6879_ (.I(_2279_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6880_ (.I(_1415_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6881_ (.I(_2281_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6882_ (.I(_2282_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6883_ (.A1(_3995_),
    .A2(_2221_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6884_ (.A1(_2280_),
    .A2(_2283_),
    .B(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6885_ (.A1(net24),
    .A2(_2278_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6886_ (.A1(_2278_),
    .A2(_2285_),
    .B(_2286_),
    .C(_1438_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6887_ (.I(_1284_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6888_ (.A1(_1412_),
    .A2(_1599_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6889_ (.A1(_1281_),
    .A2(_1250_),
    .A3(_2287_),
    .A4(_2288_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6890_ (.A1(net22),
    .A2(_2289_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6891_ (.A1(_3946_),
    .A2(_2289_),
    .B(_2290_),
    .C(_1438_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6892_ (.A1(_1283_),
    .A2(_1309_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6893_ (.I(_2291_),
    .Z(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6894_ (.I(_1091_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6895_ (.A1(_2293_),
    .A2(_1274_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6896_ (.A1(_3972_),
    .A2(_1286_),
    .B(_1577_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6897_ (.A1(_1262_),
    .A2(_2292_),
    .B1(_2294_),
    .B2(_2295_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6898_ (.I(_2281_),
    .Z(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6899_ (.A1(_1570_),
    .A2(_1259_),
    .A3(_1602_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6900_ (.I(_1611_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6901_ (.I(_2299_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6902_ (.I(_1255_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6903_ (.I(_2301_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6904_ (.A1(_2297_),
    .A2(_1276_),
    .B1(_2292_),
    .B2(_2298_),
    .C1(_2300_),
    .C2(_2302_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6905_ (.A1(_1421_),
    .A2(_2296_),
    .A3(_2303_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6906_ (.A1(net23),
    .A2(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6907_ (.A1(_3931_),
    .A2(_2304_),
    .B(_2305_),
    .C(_1635_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6908_ (.A1(_0638_),
    .A2(_0661_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6909_ (.A1(_3900_),
    .A2(_3997_),
    .A3(_4076_),
    .A4(_4267_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6910_ (.A1(_0359_),
    .A2(_0433_),
    .A3(_0564_),
    .A4(_2307_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6911_ (.A1(_2306_),
    .A2(_0733_),
    .A3(_2308_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6912_ (.A1(_0878_),
    .A2(_2309_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6913_ (.A1(_2226_),
    .A2(_2310_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6914_ (.I(_1613_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6915_ (.I(_1371_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6916_ (.A1(_1103_),
    .A2(_1072_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6917_ (.A1(_2313_),
    .A2(_1605_),
    .A3(_2314_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6918_ (.A1(_1239_),
    .A2(_2312_),
    .A3(_1598_),
    .A4(_2315_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6919_ (.A1(_1291_),
    .A2(_1598_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6920_ (.A1(_2316_),
    .A2(_2317_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6921_ (.I(_3902_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6922_ (.A1(_1251_),
    .A2(_1401_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6923_ (.A1(_4194_),
    .A2(_1398_),
    .A3(_1399_),
    .B(_2320_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6924_ (.A1(_2226_),
    .A2(_2321_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6925_ (.I(_1645_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6926_ (.A1(_2323_),
    .A2(_0896_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6927_ (.A1(_4009_),
    .A2(_1588_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6928_ (.A1(_0436_),
    .A2(_1386_),
    .B(_2325_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6929_ (.A1(_2319_),
    .A2(_2322_),
    .A3(_2324_),
    .A4(_2326_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6930_ (.A1(_1575_),
    .A2(_1373_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6931_ (.A1(_4008_),
    .A2(_1408_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6932_ (.A1(_4006_),
    .A2(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6933_ (.A1(_1732_),
    .A2(_2330_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6934_ (.A1(_4121_),
    .A2(_2291_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6935_ (.A1(_2328_),
    .A2(_2331_),
    .B(_2332_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6936_ (.A1(_1392_),
    .A2(_2333_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6937_ (.A1(_2311_),
    .A2(_2318_),
    .A3(_2327_),
    .A4(_2334_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6938_ (.A1(_1324_),
    .A2(_2312_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6939_ (.I(_1713_),
    .Z(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6940_ (.A1(_1647_),
    .A2(_1581_),
    .A3(_2337_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6941_ (.A1(_2336_),
    .A2(_2338_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6942_ (.I(_1317_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6943_ (.A1(_1298_),
    .A2(_2222_),
    .B(_1609_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6944_ (.I(_2314_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6945_ (.A1(_0495_),
    .A2(_2342_),
    .B(_1606_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6946_ (.I(_1376_),
    .Z(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6947_ (.I(_2344_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6948_ (.A1(_2345_),
    .A2(_2231_),
    .A3(_2239_),
    .A4(_2292_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6949_ (.A1(_2341_),
    .A2(_2343_),
    .A3(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6950_ (.A1(_2281_),
    .A2(_1276_),
    .B(_1248_),
    .C(_2159_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6951_ (.A1(_1306_),
    .A2(_2296_),
    .A3(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6952_ (.A1(_1613_),
    .A2(_1595_),
    .B(_1065_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6953_ (.A1(_2340_),
    .A2(_2347_),
    .A3(_2349_),
    .A4(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6954_ (.A1(_2335_),
    .A2(_2339_),
    .A3(_2351_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6955_ (.I(_2300_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6956_ (.I(_1556_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6957_ (.I(_2354_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6958_ (.I(_3950_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6959_ (.A1(_3913_),
    .A2(_1288_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6960_ (.A1(_1327_),
    .A2(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6961_ (.A1(_2356_),
    .A2(_2358_),
    .B(net26),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6962_ (.I(_2220_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6963_ (.I(_2360_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6964_ (.I(_2361_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6965_ (.A1(_2362_),
    .A2(_1264_),
    .A3(_2358_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6966_ (.A1(_2355_),
    .A2(_2359_),
    .A3(_2363_),
    .B1(_1577_),
    .B2(_2275_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6967_ (.A1(_2353_),
    .A2(_2364_),
    .B(_2352_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6968_ (.A1(net49),
    .A2(_2352_),
    .B(_2365_),
    .C(_1438_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6969_ (.I(net25),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6970_ (.A1(_2283_),
    .A2(_1276_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6971_ (.I(_2332_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6972_ (.A1(_1082_),
    .A2(_1263_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6973_ (.A1(_1107_),
    .A2(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6974_ (.A1(_1394_),
    .A2(_2370_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6975_ (.A1(_3932_),
    .A2(_3985_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6976_ (.A1(_1267_),
    .A2(_2360_),
    .A3(_2236_),
    .A4(_2372_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6977_ (.A1(_2368_),
    .A2(_2371_),
    .A3(_2373_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6978_ (.I(_1687_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6979_ (.I(_2273_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6980_ (.I(_1107_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6981_ (.A1(_1728_),
    .A2(_1415_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6982_ (.I(_2378_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6983_ (.A1(_2375_),
    .A2(_2376_),
    .A3(_2377_),
    .A4(_2379_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6984_ (.I(_1609_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6985_ (.A1(_1286_),
    .A2(_2235_),
    .A3(_3985_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6986_ (.I(_1087_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6987_ (.A1(_1573_),
    .A2(_2382_),
    .B(_2383_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6988_ (.A1(_2159_),
    .A2(_1075_),
    .A3(_2381_),
    .A4(_2384_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6989_ (.A1(_2343_),
    .A2(_2385_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6990_ (.A1(_2374_),
    .A2(_2380_),
    .A3(_2386_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6991_ (.A1(_2296_),
    .A2(_2367_),
    .A3(_2335_),
    .A4(_2387_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6992_ (.I(_1735_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6993_ (.I(_1090_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6994_ (.I(_2390_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6995_ (.I(_2370_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6996_ (.A1(_2391_),
    .A2(_1087_),
    .B(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6997_ (.A1(_1327_),
    .A2(_2393_),
    .B(_1100_),
    .C(_4279_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6998_ (.A1(_1258_),
    .A2(_2272_),
    .B(_2394_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6999_ (.A1(_2366_),
    .A2(_2282_),
    .A3(_2395_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7000_ (.I(_1556_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7001_ (.I(_2397_),
    .Z(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7002_ (.A1(_1741_),
    .A2(_2389_),
    .B(_2396_),
    .C(_2398_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7003_ (.I(_2299_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7004_ (.A1(_1718_),
    .A2(_2399_),
    .B(_2400_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7005_ (.I(_1632_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7006_ (.A1(_2388_),
    .A2(_2401_),
    .B(_2402_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7007_ (.A1(_2366_),
    .A2(_2388_),
    .B(_2403_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7008_ (.I(_1303_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7009_ (.A1(_1288_),
    .A2(_2404_),
    .A3(_2291_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7010_ (.A1(_2218_),
    .A2(_2222_),
    .A3(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7011_ (.I(_1304_),
    .Z(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7012_ (.I(_2407_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7013_ (.A1(_2319_),
    .A2(_3972_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7014_ (.A1(_2375_),
    .A2(_2282_),
    .B(_2409_),
    .C(_3932_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7015_ (.A1(_1570_),
    .A2(_2408_),
    .B(_2368_),
    .C(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7016_ (.A1(_2340_),
    .A2(_2406_),
    .A3(_2411_),
    .Z(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7017_ (.A1(_2263_),
    .A2(_2400_),
    .B(_2412_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7018_ (.I(_4187_),
    .Z(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7019_ (.I(_2414_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7020_ (.A1(_3977_),
    .A2(_2412_),
    .B(_2413_),
    .C(_2415_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7021_ (.A1(_2265_),
    .A2(_2400_),
    .B(_2412_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7022_ (.A1(_3976_),
    .A2(_2412_),
    .B(_2416_),
    .C(_2415_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7023_ (.A1(_1645_),
    .A2(_1503_),
    .A3(_1625_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7024_ (.A1(_3906_),
    .A2(_1612_),
    .A3(_2417_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7025_ (.A1(_1573_),
    .A2(_1616_),
    .B1(_1617_),
    .B2(_3951_),
    .C(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7026_ (.A1(_1600_),
    .A2(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7027_ (.I(_2420_),
    .Z(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7028_ (.I(_2421_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7029_ (.I(_2420_),
    .Z(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7030_ (.I(_1385_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7031_ (.A1(_4215_),
    .A2(_2424_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7032_ (.A1(_1673_),
    .A2(_2398_),
    .B(_2425_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7033_ (.A1(_2423_),
    .A2(_2426_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7034_ (.A1(_4138_),
    .A2(_2422_),
    .B(_2427_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7035_ (.I(_1272_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7036_ (.A1(_1531_),
    .A2(_2428_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7037_ (.A1(_0310_),
    .A2(_2397_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7038_ (.A1(_1600_),
    .A2(_2419_),
    .A3(_2429_),
    .A4(_2430_),
    .Z(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7039_ (.A1(_4293_),
    .A2(_2422_),
    .B(_2431_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7040_ (.A1(_0992_),
    .A2(_2398_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7041_ (.I(_2428_),
    .Z(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7042_ (.A1(_1532_),
    .A2(_2433_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7043_ (.A1(_1600_),
    .A2(_2419_),
    .A3(_2432_),
    .A4(_2434_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7044_ (.A1(_0320_),
    .A2(_2422_),
    .B(_2435_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7045_ (.I(_2345_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7046_ (.I(_2376_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7047_ (.A1(_1344_),
    .A2(_2437_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7048_ (.A1(_2258_),
    .A2(_2436_),
    .B(_2438_),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7049_ (.A1(_0462_),
    .A2(_2423_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7050_ (.A1(_2422_),
    .A2(_2439_),
    .B(_2440_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7051_ (.I(_2424_),
    .Z(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7052_ (.I(_2424_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7053_ (.A1(_1350_),
    .A2(_2442_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7054_ (.A1(_1660_),
    .A2(_2441_),
    .B(_2443_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7055_ (.I0(_2444_),
    .I1(_0516_),
    .S(_2421_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7056_ (.I(_2445_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7057_ (.A1(_2063_),
    .A2(_2376_),
    .B(_1426_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7058_ (.I0(_2446_),
    .I1(_0627_),
    .S(_2421_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7059_ (.I(_2447_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7060_ (.A1(_1167_),
    .A2(_2433_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7061_ (.A1(_0730_),
    .A2(_2436_),
    .B(_2448_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7062_ (.I0(_2449_),
    .I1(_0753_),
    .S(_2421_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7063_ (.I(_2450_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7064_ (.I0(_1176_),
    .I1(_2267_),
    .S(_2436_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7065_ (.A1(_0856_),
    .A2(_2423_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7066_ (.A1(_2423_),
    .A2(_2451_),
    .B(_2452_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7067_ (.I(_1437_),
    .Z(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7068_ (.A1(_2453_),
    .A2(_1607_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7069_ (.I(_1281_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7070_ (.I(_2454_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7071_ (.I(_3955_),
    .Z(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7072_ (.I(_2456_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7073_ (.A1(_2455_),
    .A2(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7074_ (.I(_2375_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7075_ (.I(_2293_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7076_ (.I(_1090_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7077_ (.I(_2461_),
    .Z(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7078_ (.A1(_2456_),
    .A2(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7079_ (.A1(_2268_),
    .A2(_2460_),
    .B1(_2372_),
    .B2(_2463_),
    .C(_2383_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7080_ (.A1(_1271_),
    .A2(_2310_),
    .A3(_2321_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7081_ (.I(_2220_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7082_ (.I(_2466_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7083_ (.A1(_2428_),
    .A2(_2463_),
    .B(_2465_),
    .C(_2467_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7084_ (.A1(_2464_),
    .A2(_2468_),
    .B(_2392_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7085_ (.I(_1413_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7086_ (.I(_2228_),
    .Z(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7087_ (.A1(_2457_),
    .A2(_1385_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7088_ (.A1(_0439_),
    .A2(_1546_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7089_ (.A1(_3913_),
    .A2(_1370_),
    .A3(_2473_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7090_ (.A1(_1377_),
    .A2(_1382_),
    .A3(_2474_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7091_ (.A1(_2471_),
    .A2(_2272_),
    .B1(_2472_),
    .B2(_2475_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7092_ (.A1(_1402_),
    .A2(_2472_),
    .B(_1593_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7093_ (.A1(_2470_),
    .A2(_2476_),
    .A3(_2477_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7094_ (.A1(_2469_),
    .A2(_2478_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7095_ (.A1(_2457_),
    .A2(_1736_),
    .B1(_2479_),
    .B2(_2292_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7096_ (.I(_2462_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7097_ (.A1(_2457_),
    .A2(_4118_),
    .B(_2481_),
    .C(_2376_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7098_ (.A1(_1302_),
    .A2(_2404_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7099_ (.I(_2483_),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7100_ (.A1(_1544_),
    .A2(_3950_),
    .B(_2484_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7101_ (.I(_1321_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7102_ (.A1(_2268_),
    .A2(_2486_),
    .B1(_3950_),
    .B2(_3916_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7103_ (.A1(_2482_),
    .A2(_2485_),
    .A3(_2487_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7104_ (.A1(_1728_),
    .A2(_2342_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7105_ (.A1(_1614_),
    .A2(_2488_),
    .A3(_2489_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7106_ (.A1(_2459_),
    .A2(_2480_),
    .B(_2490_),
    .C(_1421_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7107_ (.I(_1437_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7108_ (.A1(_2458_),
    .A2(_2491_),
    .B(_2492_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7109_ (.I(_2414_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7110_ (.A1(_1687_),
    .A2(_1284_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7111_ (.I(_2494_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7112_ (.I(_2495_),
    .Z(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7113_ (.I(_1085_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7114_ (.I(_2497_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7115_ (.A1(_2310_),
    .A2(_2321_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7116_ (.A1(_1270_),
    .A2(_2499_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7117_ (.I(_2500_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7118_ (.I(_2501_),
    .Z(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7119_ (.A1(_2357_),
    .A2(_2498_),
    .A3(_2502_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7120_ (.I(_2301_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7121_ (.I(_2229_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7122_ (.A1(_2504_),
    .A2(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7123_ (.A1(_2377_),
    .A2(_2372_),
    .B(_2503_),
    .C(_2506_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7124_ (.A1(_1425_),
    .A2(_1401_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7125_ (.A1(_2288_),
    .A2(_2475_),
    .A3(_2508_),
    .B1(_2235_),
    .B2(_3931_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7126_ (.A1(_2507_),
    .A2(_2509_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7127_ (.A1(_3931_),
    .A2(_2235_),
    .B(_2487_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7128_ (.A1(_2408_),
    .A2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7129_ (.A1(_1431_),
    .A2(_1099_),
    .A3(_2485_),
    .A4(_2512_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7130_ (.A1(_2489_),
    .A2(_2513_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7131_ (.I(_1298_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7132_ (.A1(_2496_),
    .A2(_2510_),
    .B1(_2514_),
    .B2(_2515_),
    .C(_2454_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7133_ (.A1(_2455_),
    .A2(_3930_),
    .B(_2493_),
    .C(_2516_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7134_ (.A1(_1096_),
    .A2(_2456_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7135_ (.A1(_3984_),
    .A2(_2517_),
    .Z(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7136_ (.A1(_1269_),
    .A2(_2518_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7137_ (.A1(_2356_),
    .A2(_2315_),
    .A3(_1626_),
    .B(_2519_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7138_ (.I(_1312_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7139_ (.A1(_2272_),
    .A2(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7140_ (.I(_1373_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7141_ (.A1(_1573_),
    .A2(_2523_),
    .B(_2518_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7142_ (.A1(_2522_),
    .A2(_2524_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7143_ (.A1(_1244_),
    .A2(_1425_),
    .B(_2525_),
    .C(_2470_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7144_ (.I(_1255_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7145_ (.I(_2527_),
    .Z(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7146_ (.I(_1734_),
    .Z(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7147_ (.I(_2372_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7148_ (.A1(_1093_),
    .A2(_1089_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7149_ (.A1(_2530_),
    .A2(_2519_),
    .B(_2531_),
    .C(_2362_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7150_ (.I(_2383_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7151_ (.A1(_2282_),
    .A2(_2519_),
    .B(_2379_),
    .C(_2533_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7152_ (.A1(_3986_),
    .A2(_2529_),
    .B1(_2532_),
    .B2(_2534_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7153_ (.A1(_2528_),
    .A2(_2535_),
    .B(_1688_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7154_ (.A1(_2459_),
    .A2(_2520_),
    .B1(_2526_),
    .B2(_2536_),
    .C(_2454_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7155_ (.A1(_2455_),
    .A2(_3984_),
    .B(_2493_),
    .C(_2537_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7156_ (.I(_2319_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7157_ (.A1(_1285_),
    .A2(\as2650.cycle[2] ),
    .A3(_1096_),
    .A4(_2456_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7158_ (.I(_1285_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7159_ (.A1(_3984_),
    .A2(_2517_),
    .B(_2540_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7160_ (.A1(_2539_),
    .A2(_2541_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7161_ (.A1(_3916_),
    .A2(_2356_),
    .A3(_1242_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7162_ (.I(_2484_),
    .Z(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7163_ (.A1(_2267_),
    .A2(_2356_),
    .A3(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7164_ (.A1(_2542_),
    .A2(_2543_),
    .A3(_2545_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7165_ (.I(_1269_),
    .Z(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7166_ (.A1(_2547_),
    .A2(_1099_),
    .B(_2377_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7167_ (.A1(_1741_),
    .A2(_2283_),
    .A3(_2389_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7168_ (.A1(_2377_),
    .A2(_2531_),
    .B1(_2542_),
    .B2(_2548_),
    .C(_2549_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7169_ (.A1(_2358_),
    .A2(_2546_),
    .B1(_2550_),
    .B2(_2280_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7170_ (.A1(_1285_),
    .A2(_1633_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7171_ (.A1(_2538_),
    .A2(_2551_),
    .B1(_2552_),
    .B2(_4037_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7172_ (.I(\as2650.cycle[4] ),
    .Z(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7173_ (.A1(_1281_),
    .A2(_2539_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7174_ (.A1(_2553_),
    .A2(_2554_),
    .B(_2402_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7175_ (.A1(_2553_),
    .A2(_2554_),
    .B(_2555_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7176_ (.A1(_2553_),
    .A2(_2554_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7177_ (.A1(\as2650.cycle[5] ),
    .A2(_2556_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7178_ (.A1(_2453_),
    .A2(_2557_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7179_ (.I(_1302_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7180_ (.A1(_2558_),
    .A2(_1635_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7181_ (.A1(\as2650.cycle[5] ),
    .A2(_2553_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7182_ (.A1(_2539_),
    .A2(_2560_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7183_ (.A1(_2558_),
    .A2(_2561_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7184_ (.A1(_2442_),
    .A2(_3916_),
    .B(_2515_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7185_ (.I(_2486_),
    .Z(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7186_ (.A1(_2268_),
    .A2(_2564_),
    .B(_1305_),
    .C(_2424_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7187_ (.I(_1298_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7188_ (.A1(_2437_),
    .A2(_2369_),
    .B(_2565_),
    .C(_2566_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7189_ (.A1(_2562_),
    .A2(_2563_),
    .B(_2567_),
    .C(_2455_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7190_ (.A1(_4037_),
    .A2(_2559_),
    .B(_2568_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7191_ (.I(_2486_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7192_ (.I(_2569_),
    .Z(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7193_ (.A1(_2355_),
    .A2(_2570_),
    .A3(_2544_),
    .B(_2515_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7194_ (.A1(_2558_),
    .A2(_2561_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7195_ (.A1(_1240_),
    .A2(_2572_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7196_ (.A1(_4010_),
    .A2(_2515_),
    .B1(_2571_),
    .B2(_2573_),
    .C(_2454_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7197_ (.A1(_2538_),
    .A2(_1240_),
    .B(_1633_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7198_ (.A1(_2574_),
    .A2(_2575_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7199_ (.I(_1432_),
    .Z(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7200_ (.A1(_1301_),
    .A2(_2576_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7201_ (.A1(\as2650.psu[7] ),
    .A2(_2267_),
    .B(_2577_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7202_ (.A1(_1176_),
    .A2(_2381_),
    .B1(_1582_),
    .B2(_2578_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7203_ (.A1(net4),
    .A2(_2381_),
    .A3(_1582_),
    .B(_2579_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7204_ (.I(_3903_),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7205_ (.I(_2581_),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7206_ (.A1(\as2650.psu[7] ),
    .A2(_2538_),
    .B(_2582_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7207_ (.A1(_2538_),
    .A2(_2580_),
    .B(_2583_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7208_ (.A1(_1599_),
    .A2(_0896_),
    .B1(_2342_),
    .B2(_0495_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7209_ (.A1(_3995_),
    .A2(_1099_),
    .B(_1604_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7210_ (.A1(_1612_),
    .A2(_2326_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7211_ (.A1(_1611_),
    .A2(_2585_),
    .B(_2586_),
    .C(_1608_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7212_ (.A1(_2584_),
    .A2(_2587_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7213_ (.A1(_2334_),
    .A2(_2350_),
    .A3(_2588_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7214_ (.A1(_1714_),
    .A2(_2234_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7215_ (.A1(_1575_),
    .A2(_2274_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7216_ (.A1(_2591_),
    .A2(_2332_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7217_ (.A1(_2158_),
    .A2(_1609_),
    .A3(_2590_),
    .A4(_2592_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7218_ (.A1(_2221_),
    .A2(_2531_),
    .B(_1106_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7219_ (.A1(_4122_),
    .A2(_2594_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7220_ (.A1(_2320_),
    .A2(_2489_),
    .B(_2593_),
    .C(_2595_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7221_ (.A1(_2236_),
    .A2(_2531_),
    .B(_1086_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7222_ (.A1(_1575_),
    .A2(_1592_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7223_ (.A1(_1291_),
    .A2(_2598_),
    .A3(_1613_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _7224_ (.A1(_3988_),
    .A2(_2284_),
    .A3(_2597_),
    .A4(_2599_),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7225_ (.A1(_1267_),
    .A2(_1287_),
    .A3(_1731_),
    .A4(_2330_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7226_ (.A1(_1313_),
    .A2(_2405_),
    .B1(_2601_),
    .B2(_2368_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7227_ (.A1(_2374_),
    .A2(_2596_),
    .A3(_2600_),
    .A4(_2602_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7228_ (.A1(_2316_),
    .A2(_2317_),
    .A3(_2589_),
    .A4(_2603_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7229_ (.I(_2604_),
    .Z(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7230_ (.I(_2605_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7231_ (.I(_2606_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7232_ (.I(_2604_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7233_ (.I(_1117_),
    .Z(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7234_ (.A1(_2219_),
    .A2(_1733_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7235_ (.I(_2610_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7236_ (.A1(_1117_),
    .A2(_4069_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7237_ (.A1(_0437_),
    .A2(_1713_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7238_ (.I(_2613_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7239_ (.A1(_2612_),
    .A2(_2614_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7240_ (.A1(_2609_),
    .A2(_2611_),
    .B(_2615_),
    .C(_2527_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7241_ (.A1(_2466_),
    .A2(_2329_),
    .B(_2465_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7242_ (.I(_2617_),
    .Z(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7243_ (.I(_2618_),
    .Z(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7244_ (.I(_2494_),
    .Z(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7245_ (.I(_2620_),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7246_ (.A1(_2616_),
    .A2(_2619_),
    .B(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7247_ (.I(_2270_),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7248_ (.A1(_2609_),
    .A2(_1729_),
    .Z(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7249_ (.A1(_2344_),
    .A2(_2466_),
    .A3(_2499_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7250_ (.A1(_2461_),
    .A2(_4046_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7251_ (.A1(_1673_),
    .A2(_2626_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7252_ (.A1(_2360_),
    .A2(_1395_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7253_ (.I(_2337_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7254_ (.I(\as2650.addr_buff[0] ),
    .Z(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7255_ (.A1(_2630_),
    .A2(_2293_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7256_ (.I(_4070_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7257_ (.I(_1094_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7258_ (.I(_2633_),
    .Z(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7259_ (.I(_1581_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7260_ (.A1(_2632_),
    .A2(_2634_),
    .B(_2635_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7261_ (.A1(_1117_),
    .A2(_1728_),
    .A3(_2239_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7262_ (.A1(_1591_),
    .A2(_2361_),
    .B1(_2612_),
    .B2(_1729_),
    .C(_2637_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7263_ (.A1(_2631_),
    .A2(_2636_),
    .B(_1430_),
    .C(_2638_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7264_ (.A1(_2627_),
    .A2(_2628_),
    .B(_2629_),
    .C(_2639_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7265_ (.A1(_2624_),
    .A2(_2625_),
    .B(_2640_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7266_ (.A1(_0917_),
    .A2(_0924_),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7267_ (.I(_2642_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7268_ (.I(_2643_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7269_ (.I(_0944_),
    .Z(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7270_ (.A1(_2645_),
    .A2(\as2650.stack[5][0] ),
    .B1(\as2650.stack[4][0] ),
    .B2(_1008_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7271_ (.A1(_2644_),
    .A2(_2646_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7272_ (.I(\as2650.psu[2] ),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7273_ (.A1(_2648_),
    .A2(\as2650.stack[7][0] ),
    .B1(\as2650.stack[6][0] ),
    .B2(_0918_),
    .C(_0953_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _7274_ (.I0(\as2650.stack[3][0] ),
    .I1(\as2650.stack[0][0] ),
    .I2(\as2650.stack[1][0] ),
    .I3(\as2650.stack[2][0] ),
    .S0(_0915_),
    .S1(_0916_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7275_ (.A1(_0976_),
    .A2(_2650_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7276_ (.A1(_2647_),
    .A2(_2649_),
    .B(_2651_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7277_ (.I(_2598_),
    .Z(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7278_ (.I(_2653_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _7279_ (.A1(_1119_),
    .A2(_2623_),
    .B1(_2616_),
    .B2(_2641_),
    .C1(_2652_),
    .C2(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7280_ (.I(_2495_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7281_ (.A1(_2609_),
    .A2(_2622_),
    .B1(_2655_),
    .B2(_2656_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7282_ (.A1(_2608_),
    .A2(_2657_),
    .B(_2582_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7283_ (.A1(_1119_),
    .A2(_2607_),
    .B(_2658_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7284_ (.I(_2606_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7285_ (.A1(_1278_),
    .A2(_1611_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7286_ (.I(_2660_),
    .Z(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7287_ (.A1(_1129_),
    .A2(_1116_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7288_ (.I(_2662_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7289_ (.I(_2660_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7290_ (.I(_1594_),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7291_ (.I(_1429_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7292_ (.A1(_2666_),
    .A2(_2629_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7293_ (.A1(\as2650.pc[0] ),
    .A2(net5),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7294_ (.I(_1128_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7295_ (.A1(_2669_),
    .A2(_4270_),
    .Z(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7296_ (.A1(_2668_),
    .A2(_2670_),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7297_ (.A1(_2667_),
    .A2(_2662_),
    .B1(_2671_),
    .B2(_2614_),
    .C(_1414_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7298_ (.A1(_1116_),
    .A2(\as2650.ins_reg[2] ),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7299_ (.A1(_2669_),
    .A2(_2673_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7300_ (.A1(_2313_),
    .A2(_1409_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7301_ (.I(_4205_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7302_ (.A1(_2675_),
    .A2(_2662_),
    .B1(_2671_),
    .B2(_2676_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7303_ (.I(_1409_),
    .Z(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7304_ (.I(_1089_),
    .Z(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7305_ (.A1(_4271_),
    .A2(_2679_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7306_ (.I(\as2650.addr_buff[1] ),
    .Z(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7307_ (.A1(_2681_),
    .A2(_2227_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7308_ (.A1(_2678_),
    .A2(_1086_),
    .A3(_2680_),
    .A4(_2682_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7309_ (.A1(net5),
    .A2(_4046_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7310_ (.A1(net6),
    .A2(_4082_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7311_ (.A1(_2684_),
    .A2(_2685_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7312_ (.A1(_2684_),
    .A2(_2685_),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7313_ (.A1(_1091_),
    .A2(_2686_),
    .A3(_2687_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7314_ (.A1(_4271_),
    .A2(_2633_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7315_ (.A1(_2678_),
    .A2(_2360_),
    .A3(_2688_),
    .A4(_2689_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7316_ (.A1(_2361_),
    .A2(_2677_),
    .B(_2683_),
    .C(_2690_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7317_ (.A1(_2625_),
    .A2(_2674_),
    .B1(_2691_),
    .B2(_1430_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7318_ (.A1(_2617_),
    .A2(_2663_),
    .B(_2692_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7319_ (.A1(_2505_),
    .A2(_2693_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7320_ (.I(_2643_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7321_ (.A1(_1037_),
    .A2(\as2650.stack[5][1] ),
    .B1(\as2650.stack[4][1] ),
    .B2(_1009_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7322_ (.A1(_2695_),
    .A2(_2696_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7323_ (.A1(_0950_),
    .A2(\as2650.stack[7][1] ),
    .B1(\as2650.stack[6][1] ),
    .B2(_0939_),
    .C(_0972_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7324_ (.I(_2698_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7325_ (.A1(\as2650.stack[3][1] ),
    .A2(_0934_),
    .B(_0937_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7326_ (.I0(\as2650.stack[1][1] ),
    .I1(\as2650.stack[0][1] ),
    .S(_0928_),
    .Z(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7327_ (.A1(\as2650.stack[2][1] ),
    .A2(_0919_),
    .B1(_0927_),
    .B2(_2701_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7328_ (.A1(_2700_),
    .A2(_2702_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7329_ (.A1(_2697_),
    .A2(_2699_),
    .B(_2703_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7330_ (.A1(_2654_),
    .A2(_2704_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7331_ (.A1(_2665_),
    .A2(_2663_),
    .B1(_2672_),
    .B2(_2694_),
    .C(_2705_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7332_ (.A1(_2664_),
    .A2(_2706_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7333_ (.A1(_2661_),
    .A2(_2663_),
    .B(_2707_),
    .C(_2606_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7334_ (.A1(_1130_),
    .A2(_2659_),
    .B(_2708_),
    .C(_2415_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7335_ (.I(_2605_),
    .Z(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7336_ (.A1(_1137_),
    .A2(_1128_),
    .A3(\as2650.pc[0] ),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7337_ (.A1(_1130_),
    .A2(_1118_),
    .B(_1139_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7338_ (.A1(_2710_),
    .A2(_2711_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7339_ (.A1(\as2650.pc[1] ),
    .A2(net6),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7340_ (.A1(_1128_),
    .A2(_4268_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7341_ (.A1(_2668_),
    .A2(_2713_),
    .B(_2714_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7342_ (.A1(\as2650.pc[2] ),
    .A2(net7),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7343_ (.I(_2716_),
    .Z(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7344_ (.A1(_2715_),
    .A2(_2717_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7345_ (.A1(_1413_),
    .A2(_1556_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7346_ (.I(_2719_),
    .Z(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7347_ (.A1(_4010_),
    .A2(_2712_),
    .B1(_2718_),
    .B2(_2720_),
    .C(_2392_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7348_ (.A1(_2619_),
    .A2(_2721_),
    .B(_2621_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7349_ (.I(_2675_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7350_ (.I(_2676_),
    .Z(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7351_ (.A1(_2255_),
    .A2(_1268_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7352_ (.A1(_2256_),
    .A2(_2634_),
    .B(_2725_),
    .C(_2281_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7353_ (.A1(_2723_),
    .A2(_2712_),
    .B1(_2718_),
    .B2(_2724_),
    .C(_2726_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7354_ (.I(_2501_),
    .Z(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7355_ (.A1(_1130_),
    .A2(_2673_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7356_ (.A1(_1138_),
    .A2(_2729_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7357_ (.A1(_2728_),
    .A2(_2730_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7358_ (.A1(_2397_),
    .A2(_2727_),
    .B(_2731_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7359_ (.I(_2628_),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7360_ (.I(_1268_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7361_ (.A1(_4268_),
    .A2(_4082_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7362_ (.A1(_0351_),
    .A2(_4252_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7363_ (.I(_2736_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7364_ (.A1(_2735_),
    .A2(_2686_),
    .A3(_2737_),
    .Z(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7365_ (.A1(_2735_),
    .A2(_2686_),
    .B(_2737_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7366_ (.A1(_2734_),
    .A2(_2738_),
    .A3(_2739_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7367_ (.A1(_1954_),
    .A2(_2679_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7368_ (.A1(_2733_),
    .A2(_2740_),
    .A3(_2741_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7369_ (.I(_1734_),
    .Z(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7370_ (.A1(_2533_),
    .A2(_2732_),
    .B(_2742_),
    .C(_2743_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7371_ (.A1(\as2650.stack[3][2] ),
    .A2(_0934_),
    .B(_0937_),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7372_ (.I0(\as2650.stack[1][2] ),
    .I1(\as2650.stack[0][2] ),
    .S(_0928_),
    .Z(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7373_ (.A1(\as2650.stack[2][2] ),
    .A2(_1006_),
    .B1(_0926_),
    .B2(_2746_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7374_ (.A1(_2645_),
    .A2(\as2650.stack[5][2] ),
    .B1(\as2650.stack[4][2] ),
    .B2(_1008_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7375_ (.A1(_2644_),
    .A2(_2748_),
    .Z(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7376_ (.A1(_2648_),
    .A2(\as2650.stack[7][2] ),
    .B1(\as2650.stack[6][2] ),
    .B2(_0918_),
    .C(_0971_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7377_ (.A1(_2745_),
    .A2(_2747_),
    .B1(_2749_),
    .B2(_2750_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7378_ (.I(_2653_),
    .Z(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7379_ (.A1(_2665_),
    .A2(_2712_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7380_ (.A1(_2721_),
    .A2(_2744_),
    .B1(_2751_),
    .B2(_2752_),
    .C(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7381_ (.A1(_2712_),
    .A2(_2722_),
    .B1(_2754_),
    .B2(_2656_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7382_ (.A1(_2709_),
    .A2(_2755_),
    .B(_2582_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7383_ (.A1(_1139_),
    .A2(_2607_),
    .B(_2756_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7384_ (.I(\as2650.pc[3] ),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7385_ (.A1(_2757_),
    .A2(_2710_),
    .Z(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7386_ (.A1(\as2650.pc[3] ),
    .A2(_0423_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7387_ (.A1(\as2650.pc[3] ),
    .A2(net8),
    .Z(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7388_ (.A1(_2759_),
    .A2(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7389_ (.A1(\as2650.pc[2] ),
    .A2(_0351_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7390_ (.I(_2762_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7391_ (.A1(_2715_),
    .A2(_2717_),
    .B(_2763_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7392_ (.A1(_2761_),
    .A2(_2764_),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7393_ (.A1(_4010_),
    .A2(_2758_),
    .B1(_2765_),
    .B2(_2720_),
    .C(_2392_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7394_ (.I(_2620_),
    .Z(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7395_ (.A1(_2619_),
    .A2(_2766_),
    .B(_2767_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7396_ (.A1(_0427_),
    .A2(_2390_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7397_ (.A1(_2217_),
    .A2(_2769_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7398_ (.A1(_2259_),
    .A2(_2228_),
    .B(_2770_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7399_ (.A1(_2723_),
    .A2(_2758_),
    .B1(_2765_),
    .B2(_2724_),
    .C(_2771_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7400_ (.A1(_1144_),
    .A2(_1138_),
    .A3(_1129_),
    .A4(_2673_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7401_ (.A1(_1137_),
    .A2(_2729_),
    .B(_2757_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7402_ (.A1(_2773_),
    .A2(_2774_),
    .B(_2728_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7403_ (.A1(_2354_),
    .A2(_2772_),
    .B(_2775_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7404_ (.I(_2229_),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7405_ (.A1(_0352_),
    .A2(_4252_),
    .Z(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7406_ (.A1(_0423_),
    .A2(_0362_),
    .Z(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7407_ (.A1(_2778_),
    .A2(_2739_),
    .A3(_2779_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7408_ (.A1(_2778_),
    .A2(_2739_),
    .B(_2779_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7409_ (.A1(_2391_),
    .A2(_2781_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7410_ (.A1(_0426_),
    .A2(_2633_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7411_ (.A1(_1087_),
    .A2(_2329_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7412_ (.A1(_2780_),
    .A2(_2782_),
    .B(_2783_),
    .C(_2784_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7413_ (.A1(_2777_),
    .A2(_2785_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7414_ (.A1(_2239_),
    .A2(_2776_),
    .B(_2786_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7415_ (.I(_2642_),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7416_ (.I(_0935_),
    .Z(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7417_ (.A1(_2645_),
    .A2(\as2650.stack[5][3] ),
    .B1(\as2650.stack[4][3] ),
    .B2(_2789_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7418_ (.A1(_2788_),
    .A2(_2790_),
    .Z(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7419_ (.I(_0917_),
    .Z(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7420_ (.A1(_0949_),
    .A2(\as2650.stack[7][3] ),
    .B1(\as2650.stack[6][3] ),
    .B2(_2792_),
    .C(_0971_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7421_ (.I(_0922_),
    .Z(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7422_ (.A1(_2794_),
    .A2(\as2650.stack[1][3] ),
    .B1(\as2650.stack[0][3] ),
    .B2(_2789_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7423_ (.A1(_2788_),
    .A2(_2795_),
    .Z(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7424_ (.I(_0925_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7425_ (.A1(\as2650.stack[2][3] ),
    .A2(_0918_),
    .B1(_2797_),
    .B2(\as2650.stack[3][3] ),
    .C(_0975_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7426_ (.A1(_2791_),
    .A2(_2793_),
    .B1(_2796_),
    .B2(_2798_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7427_ (.I(_2653_),
    .Z(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7428_ (.I(_1594_),
    .Z(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7429_ (.A1(_2801_),
    .A2(_2758_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7430_ (.A1(_2766_),
    .A2(_2787_),
    .B1(_2799_),
    .B2(_2800_),
    .C(_2802_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7431_ (.A1(_2758_),
    .A2(_2768_),
    .B1(_2803_),
    .B2(_2656_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7432_ (.A1(_2709_),
    .A2(_2804_),
    .B(_2582_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7433_ (.A1(_1145_),
    .A2(_2607_),
    .B(_2805_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7434_ (.A1(_1144_),
    .A2(_2710_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7435_ (.A1(_1151_),
    .A2(_2806_),
    .Z(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7436_ (.A1(\as2650.pc[4] ),
    .A2(_0559_),
    .Z(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7437_ (.A1(_2715_),
    .A2(_2716_),
    .B(_2760_),
    .C(_2763_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7438_ (.A1(_2759_),
    .A2(_2809_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7439_ (.A1(_2808_),
    .A2(_2810_),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7440_ (.A1(_2614_),
    .A2(_2811_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7441_ (.A1(_2611_),
    .A2(_2807_),
    .B(_2812_),
    .C(_2302_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7442_ (.A1(_2619_),
    .A2(_2813_),
    .B(_2767_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7443_ (.A1(_1152_),
    .A2(_2773_),
    .Z(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7444_ (.A1(_2313_),
    .A2(_1591_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7445_ (.I(\as2650.addr_buff[4] ),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7446_ (.I(_1095_),
    .Z(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7447_ (.A1(_2031_),
    .A2(_2818_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7448_ (.A1(_2817_),
    .A2(_2521_),
    .B1(_2675_),
    .B2(_2807_),
    .C(_2819_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7449_ (.A1(_2816_),
    .A2(_2811_),
    .B(_2820_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7450_ (.A1(_2728_),
    .A2(_2815_),
    .B1(_2821_),
    .B2(_2345_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7451_ (.A1(_2498_),
    .A2(_2822_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7452_ (.I(_0423_),
    .Z(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7453_ (.A1(_2824_),
    .A2(_0362_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7454_ (.A1(_0558_),
    .A2(_0412_),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7455_ (.I(_2826_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7456_ (.A1(_2825_),
    .A2(_2781_),
    .A3(_2827_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7457_ (.I(_2634_),
    .Z(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7458_ (.A1(_2825_),
    .A2(_2781_),
    .B(_2827_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7459_ (.A1(_2829_),
    .A2(_2830_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7460_ (.A1(_2031_),
    .A2(_2227_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7461_ (.A1(_2784_),
    .A2(_2832_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7462_ (.A1(_2828_),
    .A2(_2831_),
    .B(_2833_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7463_ (.A1(_2529_),
    .A2(_2823_),
    .A3(_2834_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7464_ (.A1(_1037_),
    .A2(\as2650.stack[5][4] ),
    .B1(\as2650.stack[4][4] ),
    .B2(_0942_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7465_ (.A1(_2695_),
    .A2(_2836_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7466_ (.A1(_0950_),
    .A2(\as2650.stack[7][4] ),
    .B1(\as2650.stack[6][4] ),
    .B2(_0939_),
    .C(_0972_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7467_ (.A1(_2645_),
    .A2(\as2650.stack[1][4] ),
    .B1(\as2650.stack[0][4] ),
    .B2(_1008_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7468_ (.A1(_2644_),
    .A2(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7469_ (.A1(\as2650.stack[2][4] ),
    .A2(_0939_),
    .B1(_2797_),
    .B2(\as2650.stack[3][4] ),
    .C(_2840_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7470_ (.A1(_2837_),
    .A2(_2838_),
    .B1(_2841_),
    .B2(_0972_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7471_ (.A1(_2801_),
    .A2(_2807_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7472_ (.A1(_2813_),
    .A2(_2835_),
    .B1(_2842_),
    .B2(_2800_),
    .C(_2843_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7473_ (.I(_2495_),
    .Z(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7474_ (.A1(_2807_),
    .A2(_2814_),
    .B1(_2844_),
    .B2(_2845_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7475_ (.I(_2581_),
    .Z(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7476_ (.A1(_2709_),
    .A2(_2846_),
    .B(_2847_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7477_ (.A1(_1152_),
    .A2(_2607_),
    .B(_2848_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7478_ (.I(_2606_),
    .Z(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7479_ (.A1(_1151_),
    .A2(_1144_),
    .A3(_2710_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7480_ (.A1(_1160_),
    .A2(_2850_),
    .Z(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7481_ (.I(_2618_),
    .Z(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7482_ (.I(\as2650.pc[5] ),
    .Z(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7483_ (.A1(_2853_),
    .A2(net1),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7484_ (.A1(_1159_),
    .A2(_1652_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7485_ (.A1(_2854_),
    .A2(_2855_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7486_ (.I(\as2650.pc[4] ),
    .Z(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7487_ (.A1(_1151_),
    .A2(net9),
    .Z(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7488_ (.A1(_2759_),
    .A2(_2858_),
    .A3(_2809_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7489_ (.A1(_2857_),
    .A2(_0560_),
    .B(_2859_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7490_ (.A1(_2856_),
    .A2(_2860_),
    .Z(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7491_ (.A1(_2344_),
    .A2(_1733_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7492_ (.I(_2862_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7493_ (.A1(_2611_),
    .A2(_2851_),
    .B1(_2861_),
    .B2(_2863_),
    .C(_2504_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7494_ (.A1(_2852_),
    .A2(_2864_),
    .B(_2767_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7495_ (.A1(_0658_),
    .A2(_2461_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7496_ (.A1(_2263_),
    .A2(_2818_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7497_ (.A1(_2217_),
    .A2(_2866_),
    .A3(_2867_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7498_ (.A1(_2723_),
    .A2(_2851_),
    .B1(_2861_),
    .B2(_2724_),
    .C(_2868_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7499_ (.A1(_2853_),
    .A2(_2857_),
    .A3(_2773_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7500_ (.A1(_2857_),
    .A2(_2773_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7501_ (.A1(_1160_),
    .A2(_2871_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7502_ (.A1(_2870_),
    .A2(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7503_ (.A1(_2728_),
    .A2(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7504_ (.A1(_2397_),
    .A2(_2869_),
    .B(_2874_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7505_ (.I(_2634_),
    .Z(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7506_ (.A1(_0559_),
    .A2(_0412_),
    .Z(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7507_ (.A1(net1),
    .A2(_0577_),
    .Z(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7508_ (.A1(_2877_),
    .A2(_2830_),
    .A3(_2878_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7509_ (.A1(_2877_),
    .A2(_2830_),
    .B(_2878_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7510_ (.A1(_2391_),
    .A2(_2880_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7511_ (.A1(_2879_),
    .A2(_2881_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7512_ (.A1(_1427_),
    .A2(_2876_),
    .B(_2628_),
    .C(_2882_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7513_ (.A1(_2533_),
    .A2(_2875_),
    .B(_2883_),
    .C(_2743_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7514_ (.A1(_2794_),
    .A2(\as2650.stack[1][5] ),
    .B1(\as2650.stack[0][5] ),
    .B2(_2789_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7515_ (.A1(_2788_),
    .A2(_2885_),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7516_ (.A1(\as2650.stack[2][5] ),
    .A2(_2792_),
    .B1(_0925_),
    .B2(\as2650.stack[3][5] ),
    .C(_0975_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7517_ (.A1(_0944_),
    .A2(\as2650.stack[5][5] ),
    .B1(\as2650.stack[4][5] ),
    .B2(_0941_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7518_ (.A1(_2643_),
    .A2(_2888_),
    .Z(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7519_ (.A1(_0949_),
    .A2(\as2650.stack[7][5] ),
    .B1(\as2650.stack[6][5] ),
    .B2(_0921_),
    .C(_0952_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7520_ (.A1(_2886_),
    .A2(_2887_),
    .B1(_2889_),
    .B2(_2890_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7521_ (.A1(_2801_),
    .A2(_2851_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7522_ (.A1(_2864_),
    .A2(_2884_),
    .B1(_2891_),
    .B2(_2800_),
    .C(_2892_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7523_ (.A1(_2851_),
    .A2(_2865_),
    .B1(_2893_),
    .B2(_2845_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7524_ (.A1(_2709_),
    .A2(_2894_),
    .B(_2847_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7525_ (.A1(_1160_),
    .A2(_2849_),
    .B(_2895_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7526_ (.I(_2605_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7527_ (.A1(\as2650.pc[6] ),
    .A2(_2853_),
    .A3(_2850_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7528_ (.I(_2853_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7529_ (.A1(_2898_),
    .A2(_2850_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7530_ (.A1(_1170_),
    .A2(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7531_ (.A1(_2897_),
    .A2(_2900_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7532_ (.I(_2610_),
    .Z(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7533_ (.A1(\as2650.pc[6] ),
    .A2(_0727_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7534_ (.I(_2903_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7535_ (.A1(_2859_),
    .A2(_2856_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7536_ (.A1(\as2650.pc[4] ),
    .A2(_0558_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7537_ (.A1(_2906_),
    .A2(_2854_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7538_ (.A1(_2855_),
    .A2(_2907_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7539_ (.A1(_2905_),
    .A2(_2908_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7540_ (.A1(_2904_),
    .A2(_2909_),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7541_ (.A1(_2902_),
    .A2(_2901_),
    .B1(_2910_),
    .B2(_2862_),
    .C(_2527_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7542_ (.A1(_2852_),
    .A2(_2911_),
    .B(_2767_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7543_ (.A1(_1169_),
    .A2(_2899_),
    .Z(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7544_ (.A1(_1169_),
    .A2(_2870_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7545_ (.A1(_1170_),
    .A2(_2870_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7546_ (.I(_2500_),
    .Z(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7547_ (.A1(_2914_),
    .A2(_2915_),
    .B(_2916_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7548_ (.I(_2675_),
    .Z(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7549_ (.A1(_2265_),
    .A2(_2818_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7550_ (.A1(_1539_),
    .A2(_2390_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7551_ (.A1(_2919_),
    .A2(_2920_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7552_ (.A1(_2918_),
    .A2(_2913_),
    .B1(_2921_),
    .B2(_2635_),
    .C(_2219_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7553_ (.A1(_2816_),
    .A2(_2910_),
    .B(_2922_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7554_ (.A1(_2917_),
    .A2(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7555_ (.A1(_0656_),
    .A2(_0577_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7556_ (.A1(_0727_),
    .A2(_0669_),
    .Z(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7557_ (.I(_2926_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7558_ (.A1(_2925_),
    .A2(_2880_),
    .A3(_2927_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7559_ (.A1(_2925_),
    .A2(_2880_),
    .B(_2927_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7560_ (.A1(_2734_),
    .A2(_2929_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7561_ (.A1(_1541_),
    .A2(_2829_),
    .B1(_2928_),
    .B2(_2930_),
    .C(_2628_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7562_ (.A1(_2533_),
    .A2(_2924_),
    .B(_2931_),
    .C(_1735_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7563_ (.A1(_2794_),
    .A2(\as2650.stack[1][6] ),
    .B1(\as2650.stack[0][6] ),
    .B2(_2789_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7564_ (.A1(_2788_),
    .A2(_2933_),
    .Z(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7565_ (.A1(\as2650.stack[2][6] ),
    .A2(_2792_),
    .B1(_2797_),
    .B2(\as2650.stack[3][6] ),
    .C(_0975_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7566_ (.A1(_2794_),
    .A2(\as2650.stack[5][6] ),
    .B1(\as2650.stack[4][6] ),
    .B2(_0941_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7567_ (.A1(_2643_),
    .A2(_2936_),
    .Z(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7568_ (.A1(_0949_),
    .A2(\as2650.stack[7][6] ),
    .B1(\as2650.stack[6][6] ),
    .B2(_2792_),
    .C(_0971_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7569_ (.A1(_2934_),
    .A2(_2935_),
    .B1(_2937_),
    .B2(_2938_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _7570_ (.A1(_2623_),
    .A2(_2913_),
    .B1(_2911_),
    .B2(_2932_),
    .C1(_2939_),
    .C2(_2654_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7571_ (.A1(_2901_),
    .A2(_2912_),
    .B1(_2940_),
    .B2(_2845_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7572_ (.A1(_2896_),
    .A2(_2941_),
    .B(_2847_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7573_ (.A1(_1170_),
    .A2(_2849_),
    .B(_2942_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7574_ (.I(\as2650.pc[7] ),
    .Z(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7575_ (.A1(_2943_),
    .A2(_2897_),
    .Z(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7576_ (.I(_2613_),
    .Z(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7577_ (.I(_2945_),
    .Z(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7578_ (.A1(\as2650.pc[7] ),
    .A2(_0727_),
    .Z(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7579_ (.A1(_1168_),
    .A2(_2084_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7580_ (.A1(_2903_),
    .A2(_2909_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7581_ (.A1(_2948_),
    .A2(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7582_ (.A1(_2947_),
    .A2(_2950_),
    .Z(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7583_ (.A1(_2946_),
    .A2(_2951_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7584_ (.A1(_2611_),
    .A2(_2944_),
    .B(_2952_),
    .C(_2302_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7585_ (.I(_2620_),
    .Z(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7586_ (.A1(_2852_),
    .A2(_2953_),
    .B(_2954_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7587_ (.A1(_2083_),
    .A2(_0669_),
    .Z(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7588_ (.A1(net3),
    .A2(_4101_),
    .Z(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7589_ (.A1(_2956_),
    .A2(_2929_),
    .B(_2957_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7590_ (.A1(_2956_),
    .A2(_2929_),
    .A3(_2957_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7591_ (.A1(_2829_),
    .A2(_2959_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7592_ (.A1(_1544_),
    .A2(_2876_),
    .B1(_2958_),
    .B2(_2960_),
    .C(_2733_),
    .ZN(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7593_ (.A1(_1177_),
    .A2(_2914_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7594_ (.A1(_0876_),
    .A2(_2390_),
    .B1(_2521_),
    .B2(_1241_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7595_ (.A1(_2378_),
    .A2(_2944_),
    .B(_2963_),
    .C(_2344_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7596_ (.A1(_2724_),
    .A2(_2951_),
    .B(_2964_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7597_ (.A1(_2502_),
    .A2(_2962_),
    .B(_2965_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7598_ (.A1(_2498_),
    .A2(_2966_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7599_ (.A1(_2529_),
    .A2(_2961_),
    .A3(_2967_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7600_ (.A1(_0945_),
    .A2(\as2650.stack[1][7] ),
    .B1(\as2650.stack[0][7] ),
    .B2(_0942_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7601_ (.A1(\as2650.stack[2][7] ),
    .A2(_1006_),
    .B1(_2797_),
    .B2(\as2650.stack[3][7] ),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7602_ (.A1(_2644_),
    .A2(_2969_),
    .B(_2970_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7603_ (.A1(_1037_),
    .A2(\as2650.stack[5][7] ),
    .B1(\as2650.stack[4][7] ),
    .B2(_0942_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7604_ (.A1(_2695_),
    .A2(_2972_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7605_ (.A1(_2648_),
    .A2(\as2650.stack[7][7] ),
    .B1(\as2650.stack[6][7] ),
    .B2(_1006_),
    .C(_0953_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7606_ (.I(_2974_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7607_ (.A1(_0976_),
    .A2(_2971_),
    .B1(_2973_),
    .B2(_2975_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7608_ (.I(_1262_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7609_ (.A1(_2665_),
    .A2(_2944_),
    .B1(_2976_),
    .B2(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7610_ (.A1(_2953_),
    .A2(_2968_),
    .B(_2978_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7611_ (.A1(_2944_),
    .A2(_2955_),
    .B1(_2979_),
    .B2(_2845_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7612_ (.A1(_2896_),
    .A2(_2980_),
    .B(_2847_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7613_ (.A1(_1177_),
    .A2(_2849_),
    .B(_2981_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7614_ (.I(_2620_),
    .Z(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7615_ (.A1(\as2650.pc[8] ),
    .A2(_1536_),
    .Z(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7616_ (.A1(_2903_),
    .A2(_2947_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7617_ (.I(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7618_ (.A1(_2943_),
    .A2(\as2650.pc[6] ),
    .B(_1536_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7619_ (.I(_2986_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7620_ (.A1(_2909_),
    .A2(_2985_),
    .B(_2987_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7621_ (.A1(_2983_),
    .A2(_2988_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7622_ (.A1(_1177_),
    .A2(_2897_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7623_ (.A1(_1188_),
    .A2(_2990_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7624_ (.I(_1255_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7625_ (.A1(_2862_),
    .A2(_2989_),
    .B1(_2991_),
    .B2(_2610_),
    .C(_2992_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7626_ (.I(_2943_),
    .Z(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7627_ (.A1(_2994_),
    .A2(_2914_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7628_ (.A1(_1189_),
    .A2(_2995_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7629_ (.A1(_2313_),
    .A2(_2989_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7630_ (.A1(_1729_),
    .A2(_2991_),
    .B(_2678_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _7631_ (.A1(_2630_),
    .A2(_2461_),
    .B1(_2997_),
    .B2(_2998_),
    .C1(_2521_),
    .C2(_2632_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7632_ (.A1(_2916_),
    .A2(_2996_),
    .B1(_2999_),
    .B2(_2666_),
    .ZN(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7633_ (.I(\as2650.addr_buff[0] ),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7634_ (.A1(_0874_),
    .A2(_4101_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7635_ (.A1(_3002_),
    .A2(_2958_),
    .B(_1095_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7636_ (.A1(_3001_),
    .A2(_3003_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7637_ (.A1(_2498_),
    .A2(_3000_),
    .B1(_3004_),
    .B2(_2733_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7638_ (.A1(_2743_),
    .A2(_3005_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7639_ (.A1(_2801_),
    .A2(_2991_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7640_ (.A1(_0956_),
    .A2(_2800_),
    .B1(_2993_),
    .B2(_3006_),
    .C(_3007_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7641_ (.I(_2617_),
    .Z(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7642_ (.A1(_3009_),
    .A2(_2993_),
    .B(_2954_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7643_ (.I(_2604_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7644_ (.A1(_2982_),
    .A2(_3008_),
    .B1(_3010_),
    .B2(_2991_),
    .C(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7645_ (.A1(_1190_),
    .A2(_2608_),
    .B(_3012_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7646_ (.A1(_2453_),
    .A2(_3013_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7647_ (.A1(_1196_),
    .A2(\as2650.pc[8] ),
    .A3(_2990_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7648_ (.A1(_1189_),
    .A2(_2990_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7649_ (.A1(_1198_),
    .A2(_3015_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7650_ (.A1(_3014_),
    .A2(_3016_),
    .ZN(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7651_ (.A1(\as2650.pc[9] ),
    .A2(_0728_),
    .Z(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7652_ (.I(_2983_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7653_ (.A1(_1188_),
    .A2(_1537_),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7654_ (.A1(_3019_),
    .A2(_2988_),
    .B(_3020_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7655_ (.A1(_3018_),
    .A2(_3021_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7656_ (.A1(_2945_),
    .A2(_3022_),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7657_ (.A1(_2902_),
    .A2(_3017_),
    .B(_3023_),
    .C(_2504_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7658_ (.A1(_2852_),
    .A2(_3024_),
    .B(_2954_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7659_ (.A1(_3001_),
    .A2(_3003_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7660_ (.A1(_2681_),
    .A2(_3026_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7661_ (.I(_1196_),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7662_ (.A1(_1188_),
    .A2(_2943_),
    .A3(_2914_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7663_ (.A1(_3028_),
    .A2(_3029_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7664_ (.A1(_1197_),
    .A2(_3015_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7665_ (.A1(_2681_),
    .A2(_1091_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7666_ (.A1(_2689_),
    .A2(_3032_),
    .B(_1415_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7667_ (.A1(_2918_),
    .A2(_3031_),
    .B1(_3022_),
    .B2(_2676_),
    .C(_3033_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7668_ (.A1(_2501_),
    .A2(_3030_),
    .B1(_3034_),
    .B2(_2666_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7669_ (.A1(_2733_),
    .A2(_3027_),
    .B1(_3035_),
    .B2(_2467_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7670_ (.A1(_2743_),
    .A2(_3036_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _7671_ (.A1(_0981_),
    .A2(_2752_),
    .B1(_3024_),
    .B2(_3037_),
    .C1(_3031_),
    .C2(_2623_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7672_ (.A1(_3017_),
    .A2(_3025_),
    .B1(_3038_),
    .B2(_2982_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7673_ (.I(_2581_),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7674_ (.A1(_2896_),
    .A2(_3039_),
    .B(_3040_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7675_ (.A1(_1198_),
    .A2(_2849_),
    .B(_3041_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7676_ (.I(\as2650.pc[10] ),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7677_ (.A1(_1204_),
    .A2(_1536_),
    .Z(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7678_ (.I(_3043_),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7679_ (.I(_3018_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7680_ (.A1(_3019_),
    .A2(_2988_),
    .A3(_3045_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7681_ (.A1(_1196_),
    .A2(_1537_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7682_ (.A1(_3020_),
    .A2(_3047_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7683_ (.A1(_3046_),
    .A2(_3048_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7684_ (.A1(_3044_),
    .A2(_3049_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7685_ (.A1(\as2650.pc[10] ),
    .A2(_3014_),
    .Z(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7686_ (.A1(_2863_),
    .A2(_3050_),
    .B1(_3051_),
    .B2(_2902_),
    .C(_2527_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7687_ (.I(_2784_),
    .Z(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7688_ (.A1(_2630_),
    .A2(_2681_),
    .A3(_3003_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7689_ (.A1(_2256_),
    .A2(_3054_),
    .Z(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7690_ (.A1(_1205_),
    .A2(_1197_),
    .A3(_3029_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7691_ (.A1(_1198_),
    .A2(_3029_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7692_ (.A1(_3042_),
    .A2(_3057_),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7693_ (.A1(_3056_),
    .A2(_3058_),
    .B(_2501_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7694_ (.A1(\as2650.addr_buff[2] ),
    .A2(_2679_),
    .Z(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7695_ (.A1(_2741_),
    .A2(_3060_),
    .Z(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7696_ (.A1(_2217_),
    .A2(_3061_),
    .B(_0438_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7697_ (.A1(_2816_),
    .A2(_3050_),
    .B1(_3051_),
    .B2(_2379_),
    .C(_3062_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7698_ (.A1(_3059_),
    .A2(_3063_),
    .B(_2467_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7699_ (.A1(_3053_),
    .A2(_3055_),
    .B(_3064_),
    .C(_1735_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7700_ (.A1(_1000_),
    .A2(_2752_),
    .B1(_3052_),
    .B2(_3065_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7701_ (.A1(_3009_),
    .A2(_3052_),
    .B(_2623_),
    .C(_2495_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7702_ (.A1(_2982_),
    .A2(_3066_),
    .B1(_3067_),
    .B2(_3051_),
    .C(_2605_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7703_ (.A1(_3042_),
    .A2(_2608_),
    .B(_3068_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7704_ (.A1(_2453_),
    .A2(_3069_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7705_ (.I(_2271_),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7706_ (.A1(_1205_),
    .A2(_3014_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7707_ (.A1(_1213_),
    .A2(_3071_),
    .Z(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7708_ (.I(_3072_),
    .Z(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7709_ (.A1(_2618_),
    .A2(_3073_),
    .B(_2777_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7710_ (.A1(\as2650.addr_buff[0] ),
    .A2(\as2650.addr_buff[1] ),
    .A3(\as2650.addr_buff[2] ),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7711_ (.A1(_3002_),
    .A2(_2958_),
    .B(_3075_),
    .C(_2227_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7712_ (.A1(\as2650.addr_buff[3] ),
    .A2(_3076_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7713_ (.A1(\as2650.addr_buff[3] ),
    .A2(_3076_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7714_ (.A1(_1396_),
    .A2(_3077_),
    .A3(_3078_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7715_ (.A1(_1212_),
    .A2(_0728_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7716_ (.A1(\as2650.pc[10] ),
    .A2(_2083_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7717_ (.A1(_3044_),
    .A2(_3049_),
    .B(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7718_ (.A1(_3080_),
    .A2(_3082_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7719_ (.A1(\as2650.addr_buff[3] ),
    .A2(_2679_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7720_ (.A1(_2783_),
    .A2(_3084_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7721_ (.A1(_1410_),
    .A2(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7722_ (.A1(_2816_),
    .A2(_3083_),
    .B1(_3072_),
    .B2(_2379_),
    .C(_3086_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7723_ (.I(\as2650.pc[11] ),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7724_ (.A1(_3088_),
    .A2(_3056_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7725_ (.A1(_2345_),
    .A2(_3087_),
    .B1(_3089_),
    .B2(_2916_),
    .C(_2467_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7726_ (.A1(_2362_),
    .A2(_3079_),
    .B(_3090_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7727_ (.A1(_2946_),
    .A2(_3083_),
    .B1(_3073_),
    .B2(_2667_),
    .C(_1414_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7728_ (.A1(_3074_),
    .A2(_3091_),
    .B(_3092_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7729_ (.A1(_1018_),
    .A2(_2977_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7730_ (.A1(_3070_),
    .A2(_3073_),
    .B(_3093_),
    .C(_3094_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7731_ (.A1(_2621_),
    .A2(_3073_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7732_ (.A1(_2496_),
    .A2(_3095_),
    .B(_3096_),
    .C(_3011_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7733_ (.A1(_1213_),
    .A2(_2659_),
    .B(_3097_),
    .C(_2415_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7734_ (.A1(_1219_),
    .A2(\as2650.pc[11] ),
    .A3(_3071_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7735_ (.A1(_1213_),
    .A2(_1205_),
    .A3(_3014_),
    .B(_1220_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7736_ (.A1(_3098_),
    .A2(_3099_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7737_ (.A1(_3043_),
    .A2(_3080_),
    .ZN(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7738_ (.A1(_3020_),
    .A2(_3047_),
    .A3(_3081_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7739_ (.A1(\as2650.pc[11] ),
    .A2(_2084_),
    .B1(_3046_),
    .B2(_3101_),
    .C(_3102_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7740_ (.A1(\as2650.pc[12] ),
    .A2(_2083_),
    .Z(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7741_ (.A1(_3103_),
    .A2(_3104_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7742_ (.A1(_2614_),
    .A2(_3105_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7743_ (.A1(_2902_),
    .A2(_3100_),
    .B(_3106_),
    .C(_2504_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7744_ (.A1(_3009_),
    .A2(_3107_),
    .B(_2954_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7745_ (.A1(_2261_),
    .A2(_3078_),
    .Z(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7746_ (.A1(_1219_),
    .A2(_3088_),
    .A3(_3056_),
    .Z(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7747_ (.A1(_3088_),
    .A2(_3056_),
    .B(_1219_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7748_ (.A1(_3110_),
    .A2(_3111_),
    .Z(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7749_ (.A1(_2676_),
    .A2(_3105_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7750_ (.I(_3100_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7751_ (.A1(_2817_),
    .A2(_1268_),
    .B(_2832_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7752_ (.A1(_2918_),
    .A2(_3114_),
    .B1(_3115_),
    .B2(_2635_),
    .C(_2219_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7753_ (.A1(_2916_),
    .A2(_3112_),
    .B1(_3113_),
    .B2(_3116_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7754_ (.A1(_2497_),
    .A2(_3117_),
    .B(_2629_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7755_ (.A1(_3053_),
    .A2(_3109_),
    .B(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _7756_ (.A1(_1031_),
    .A2(_2752_),
    .B1(_3107_),
    .B2(_3119_),
    .C1(_3114_),
    .C2(_2271_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7757_ (.A1(_3100_),
    .A2(_3108_),
    .B1(_3120_),
    .B2(_2982_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7758_ (.A1(_2896_),
    .A2(_3121_),
    .B(_3040_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7759_ (.A1(_1221_),
    .A2(_2659_),
    .B(_3122_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7760_ (.A1(_1227_),
    .A2(_3098_),
    .Z(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7761_ (.A1(_1227_),
    .A2(_3110_),
    .Z(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7762_ (.A1(_2263_),
    .A2(_2462_),
    .B1(_2918_),
    .B2(_3123_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7763_ (.A1(_2502_),
    .A2(_3124_),
    .B1(_3125_),
    .B2(_2428_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7764_ (.A1(_2817_),
    .A2(_3078_),
    .B(_2867_),
    .C(_3053_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7765_ (.A1(_2618_),
    .A2(_3123_),
    .B1(_3126_),
    .B2(_2362_),
    .C(_3127_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7766_ (.A1(_1043_),
    .A2(_2977_),
    .B1(_3123_),
    .B2(_2665_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7767_ (.A1(_2506_),
    .A2(_3128_),
    .B(_3129_),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7768_ (.A1(_1254_),
    .A2(_0437_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7769_ (.I(_2629_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7770_ (.A1(_3131_),
    .A2(_3132_),
    .B(_2621_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7771_ (.A1(_2496_),
    .A2(_3130_),
    .B1(_3133_),
    .B2(_3123_),
    .C(_3011_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7772_ (.I(_2414_),
    .Z(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7773_ (.A1(_1227_),
    .A2(_2659_),
    .B(_3134_),
    .C(_3135_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7774_ (.A1(_1226_),
    .A2(_3098_),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7775_ (.A1(_1234_),
    .A2(_3136_),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7776_ (.A1(_3132_),
    .A2(_3009_),
    .B(_3137_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7777_ (.A1(\as2650.pc[13] ),
    .A2(_3110_),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7778_ (.A1(\as2650.pc[14] ),
    .A2(_3139_),
    .B(_2497_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7779_ (.A1(\as2650.pc[14] ),
    .A2(_3139_),
    .B(_3140_),
    .C(_2502_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7780_ (.A1(_1272_),
    .A2(_2383_),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7781_ (.A1(_2265_),
    .A2(_2462_),
    .B1(_2723_),
    .B2(_3137_),
    .C(_3142_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7782_ (.A1(_3053_),
    .A2(_2919_),
    .B(_3143_),
    .C(_2946_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7783_ (.A1(_3141_),
    .A2(_3144_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7784_ (.A1(_3138_),
    .A2(_3145_),
    .B(_2528_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7785_ (.A1(_1054_),
    .A2(_2654_),
    .B1(_3137_),
    .B2(_2271_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7786_ (.A1(_2661_),
    .A2(_3147_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7787_ (.A1(_2661_),
    .A2(_3137_),
    .B1(_3146_),
    .B2(_3148_),
    .C(_3011_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7788_ (.A1(_1234_),
    .A2(_2608_),
    .B(_3149_),
    .C(_3135_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7789_ (.I(_2460_),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7790_ (.A1(_2570_),
    .A2(_4062_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7791_ (.I(_2216_),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7792_ (.I(_3152_),
    .Z(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7793_ (.A1(_3153_),
    .A2(_4131_),
    .B(_3150_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7794_ (.I(_1318_),
    .Z(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7795_ (.A1(_3150_),
    .A2(_4183_),
    .B1(_3151_),
    .B2(_3154_),
    .C(_3155_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7796_ (.I(_1258_),
    .Z(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7797_ (.I(_1566_),
    .Z(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7798_ (.I(_1563_),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7799_ (.I(_3159_),
    .Z(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7800_ (.I(_1585_),
    .Z(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7801_ (.I(_3161_),
    .Z(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7802_ (.I(_0912_),
    .Z(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7803_ (.I(_1386_),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7804_ (.A1(_1014_),
    .A2(_1387_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7805_ (.A1(_4108_),
    .A2(_3164_),
    .B(_3165_),
    .C(_0902_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7806_ (.A1(_4222_),
    .A2(_3162_),
    .B1(_3163_),
    .B2(_2652_),
    .C(_3166_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7807_ (.A1(_1564_),
    .A2(_3167_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7808_ (.I(_4029_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7809_ (.A1(_3160_),
    .A2(_1842_),
    .B(_3168_),
    .C(_3169_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7810_ (.A1(_3158_),
    .A2(_1335_),
    .B(_3170_),
    .C(_1550_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7811_ (.A1(_1717_),
    .A2(_1529_),
    .B(_3157_),
    .C(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7812_ (.A1(_0898_),
    .A2(_2316_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7813_ (.A1(_1270_),
    .A2(_1594_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7814_ (.A1(_1256_),
    .A2(_1273_),
    .A3(_2523_),
    .A4(_3174_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7815_ (.A1(_1069_),
    .A2(_1085_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7816_ (.A1(_1246_),
    .A2(_2598_),
    .A3(_2291_),
    .A4(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7817_ (.A1(_1292_),
    .A2(_1296_),
    .B(_3177_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7818_ (.A1(_1527_),
    .A2(_2288_),
    .B(_1580_),
    .C(_3178_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7819_ (.A1(_3994_),
    .A2(_1065_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7820_ (.A1(_1289_),
    .A2(_3175_),
    .A3(_3179_),
    .A4(_3180_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7821_ (.A1(_1316_),
    .A2(_1603_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7822_ (.A1(_3181_),
    .A2(_3182_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7823_ (.A1(_1271_),
    .A2(_1587_),
    .Z(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7824_ (.A1(_3998_),
    .A2(_1555_),
    .A3(_1806_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7825_ (.A1(_1104_),
    .A2(_2337_),
    .A3(_3185_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7826_ (.A1(_1324_),
    .A2(_3184_),
    .A3(_2343_),
    .A4(_3186_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7827_ (.A1(_2523_),
    .A2(_2342_),
    .B1(_1579_),
    .B2(_3962_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7828_ (.I(_4123_),
    .Z(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7829_ (.A1(_4119_),
    .A2(_3189_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7830_ (.A1(_1093_),
    .A2(_3920_),
    .ZN(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7831_ (.A1(_2216_),
    .A2(_3191_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7832_ (.A1(_1806_),
    .A2(_4118_),
    .B1(_2633_),
    .B2(_3990_),
    .C(_1304_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7833_ (.A1(_3192_),
    .A2(_3193_),
    .B(_1257_),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7834_ (.A1(_1806_),
    .A2(_3188_),
    .B1(_3190_),
    .B2(_1313_),
    .C(_3194_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7835_ (.A1(_3173_),
    .A2(_3183_),
    .A3(_3187_),
    .A4(_3195_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7836_ (.I(_3196_),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7837_ (.I(_2231_),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7838_ (.A1(_1849_),
    .A2(_3198_),
    .B1(_1622_),
    .B2(_0872_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7839_ (.A1(_3172_),
    .A2(_3197_),
    .A3(_3199_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7840_ (.A1(_3156_),
    .A2(_3200_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7841_ (.I(_3196_),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7842_ (.I(_3202_),
    .Z(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7843_ (.A1(_4216_),
    .A2(_3203_),
    .B(_1633_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7844_ (.A1(_3201_),
    .A2(_3204_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7845_ (.I(_2569_),
    .Z(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7846_ (.A1(_3205_),
    .A2(_4244_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7847_ (.I(_2471_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7848_ (.A1(_2570_),
    .A2(_4236_),
    .B(_3206_),
    .C(_3207_),
    .ZN(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7849_ (.A1(_3150_),
    .A2(_0301_),
    .B(_3155_),
    .ZN(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7850_ (.I(_1387_),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7851_ (.A1(_0978_),
    .A2(_3210_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7852_ (.A1(_1666_),
    .A2(_1388_),
    .B(_3211_),
    .C(_1389_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7853_ (.I(_1563_),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7854_ (.A1(_0308_),
    .A2(_3162_),
    .B(_3212_),
    .C(_3213_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7855_ (.A1(_2156_),
    .A2(_2704_),
    .B(_3214_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7856_ (.A1(_3160_),
    .A2(_4251_),
    .B(_1567_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7857_ (.A1(_3158_),
    .A2(_4261_),
    .B1(_3215_),
    .B2(_3216_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7858_ (.A1(_1529_),
    .A2(_3217_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7859_ (.A1(_2251_),
    .A2(_1643_),
    .B(_1577_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7860_ (.A1(_1687_),
    .A2(_2273_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7861_ (.I(_3220_),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7862_ (.A1(_4267_),
    .A2(_1721_),
    .B1(_3221_),
    .B2(_1335_),
    .C(_3202_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7863_ (.A1(_3208_),
    .A2(_3209_),
    .B1(_3218_),
    .B2(_3219_),
    .C(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7864_ (.I(_1632_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7865_ (.A1(_0965_),
    .A2(_3203_),
    .B(_3224_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7866_ (.A1(_3223_),
    .A2(_3225_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7867_ (.I(_1293_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7868_ (.A1(_3152_),
    .A2(_0393_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7869_ (.A1(_3152_),
    .A2(_0386_),
    .B(_3227_),
    .C(_2547_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7870_ (.A1(_3207_),
    .A2(_0349_),
    .B(_3226_),
    .C(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7871_ (.I(\as2650.overflow ),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7872_ (.A1(_2648_),
    .A2(_1387_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7873_ (.A1(_3230_),
    .A2(_3210_),
    .B(_3231_),
    .C(_0903_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7874_ (.A1(_0501_),
    .A2(_3162_),
    .B1(_0913_),
    .B2(_2751_),
    .C(_3232_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7875_ (.A1(_3213_),
    .A2(_3233_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7876_ (.A1(_3160_),
    .A2(_4092_),
    .B(_3234_),
    .C(_1567_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7877_ (.A1(_3158_),
    .A2(_1345_),
    .B(_3235_),
    .C(_1550_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7878_ (.A1(_1725_),
    .A2(_1529_),
    .B(_3157_),
    .C(_3236_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7879_ (.A1(_1953_),
    .A2(_3198_),
    .B1(_1623_),
    .B2(_4261_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7880_ (.A1(_3197_),
    .A2(_3229_),
    .A3(_3237_),
    .A4(_3238_),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7881_ (.I(_3196_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7882_ (.A1(_0993_),
    .A2(_3240_),
    .B(_3224_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7883_ (.A1(_3239_),
    .A2(_3241_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7884_ (.I(_1437_),
    .Z(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7885_ (.A1(_2569_),
    .A2(_0454_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7886_ (.A1(_2564_),
    .A2(_0460_),
    .B(_3243_),
    .C(_2547_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7887_ (.A1(_3207_),
    .A2(_0492_),
    .B(_3226_),
    .C(_3244_),
    .ZN(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7888_ (.I(_1533_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7889_ (.I(_1528_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7890_ (.A1(_1380_),
    .A2(_1378_),
    .A3(_0911_),
    .ZN(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7891_ (.A1(_4095_),
    .A2(_3248_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7892_ (.A1(_1651_),
    .A2(_3248_),
    .B(_3249_),
    .C(_0902_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7893_ (.A1(_1210_),
    .A2(_3161_),
    .B1(_3163_),
    .B2(_2799_),
    .C(_3250_),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7894_ (.A1(_1564_),
    .A2(_3251_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7895_ (.A1(_3213_),
    .A2(_4261_),
    .B(_3252_),
    .C(_3169_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7896_ (.A1(_3158_),
    .A2(_1351_),
    .B(_3253_),
    .C(_1550_),
    .ZN(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7897_ (.A1(_3246_),
    .A2(_3247_),
    .B(_3157_),
    .C(_3254_),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7898_ (.A1(_0433_),
    .A2(_1720_),
    .B1(_3220_),
    .B2(_1345_),
    .C(_3196_),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7899_ (.I(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7900_ (.A1(_3245_),
    .A2(_3255_),
    .A3(_3257_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7901_ (.A1(_1344_),
    .A2(_3240_),
    .B(_3258_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7902_ (.A1(_3242_),
    .A2(_3259_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7903_ (.I(_2471_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7904_ (.A1(_3153_),
    .A2(_0556_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7905_ (.A1(_2570_),
    .A2(_0594_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7906_ (.A1(_3260_),
    .A2(_3261_),
    .A3(_3262_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7907_ (.A1(_3260_),
    .A2(_0548_),
    .B(_1525_),
    .C(_3263_),
    .ZN(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7908_ (.A1(_0564_),
    .A2(_1721_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7909_ (.I(_1684_),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7910_ (.I(\as2650.psu[4] ),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7911_ (.A1(_4036_),
    .A2(_3210_),
    .B(_1389_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7912_ (.A1(_3267_),
    .A2(_1388_),
    .B(_3268_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7913_ (.A1(_0615_),
    .A2(_0896_),
    .B1(_2156_),
    .B2(_2842_),
    .C(_3269_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7914_ (.A1(_3213_),
    .A2(_0370_),
    .B(_1566_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7915_ (.A1(_3160_),
    .A2(_3270_),
    .B(_3271_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7916_ (.A1(_3266_),
    .A2(_0586_),
    .B(_3272_),
    .C(_1643_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7917_ (.I(_1258_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7918_ (.A1(_1535_),
    .A2(_3247_),
    .B(_3274_),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7919_ (.A1(_1351_),
    .A2(_3221_),
    .B1(_3273_),
    .B2(_3275_),
    .C(_3202_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7920_ (.A1(_3265_),
    .A2(_3276_),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7921_ (.A1(_1350_),
    .A2(_3240_),
    .B(_3040_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7922_ (.A1(_3264_),
    .A2(_3277_),
    .B(_3278_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7923_ (.A1(_3205_),
    .A2(_0682_),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7924_ (.A1(_3153_),
    .A2(_0654_),
    .B(_2481_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7925_ (.I(_1318_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7926_ (.A1(_3150_),
    .A2(_2062_),
    .B1(_3279_),
    .B2(_3280_),
    .C(_3281_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7927_ (.A1(_1667_),
    .A2(_3164_),
    .B(_0903_),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7928_ (.A1(\as2650.psu[5] ),
    .A2(_3210_),
    .B(_3283_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7929_ (.A1(_0574_),
    .A2(_3161_),
    .B1(_3163_),
    .B2(_2891_),
    .C(_1563_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7930_ (.A1(_3159_),
    .A2(_1351_),
    .B1(_3284_),
    .B2(_3285_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7931_ (.A1(_3169_),
    .A2(_3286_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7932_ (.A1(_1684_),
    .A2(_1361_),
    .ZN(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7933_ (.A1(_1528_),
    .A2(_3287_),
    .A3(_3288_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7934_ (.A1(_1428_),
    .A2(_3247_),
    .B(_3274_),
    .C(_3289_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7935_ (.A1(_1356_),
    .A2(_3221_),
    .B(_3202_),
    .C(_3290_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7936_ (.A1(_2306_),
    .A2(_3198_),
    .B(_3282_),
    .C(_3291_),
    .ZN(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7937_ (.A1(_1157_),
    .A2(_3240_),
    .B(_3224_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7938_ (.A1(_3292_),
    .A2(_3293_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7939_ (.A1(_3152_),
    .A2(_0726_),
    .ZN(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7940_ (.A1(_3205_),
    .A2(_0722_),
    .B(_2547_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7941_ (.I(_1524_),
    .Z(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7942_ (.A1(_3260_),
    .A2(_1518_),
    .B1(_3294_),
    .B2(_3295_),
    .C(_3296_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7943_ (.A1(_1668_),
    .A2(_3164_),
    .B(_0903_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7944_ (.A1(net27),
    .A2(_1388_),
    .B(_3298_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7945_ (.A1(_1233_),
    .A2(_3161_),
    .B1(_3163_),
    .B2(_2939_),
    .C(_3159_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7946_ (.A1(_1564_),
    .A2(_1356_),
    .B1(_3299_),
    .B2(_3300_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7947_ (.A1(_3169_),
    .A2(_3301_),
    .ZN(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7948_ (.A1(_1567_),
    .A2(_1624_),
    .B(_3302_),
    .C(_1528_),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7949_ (.A1(_1739_),
    .A2(_3247_),
    .B(_3303_),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7950_ (.A1(_0715_),
    .A2(_1623_),
    .B1(_3304_),
    .B2(_3157_),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7951_ (.A1(_0733_),
    .A2(_1721_),
    .B(_3297_),
    .C(_3305_),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7952_ (.A1(_1167_),
    .A2(_3197_),
    .B(_3040_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7953_ (.A1(_3203_),
    .A2(_3306_),
    .B(_3307_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7954_ (.A1(_3153_),
    .A2(_0886_),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7955_ (.A1(_3205_),
    .A2(_0868_),
    .B(_3207_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7956_ (.A1(_3260_),
    .A2(_0862_),
    .B1(_3308_),
    .B2(_3309_),
    .C(_1525_),
    .ZN(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7957_ (.I(\as2650.psu[7] ),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7958_ (.A1(_1636_),
    .A2(_3248_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7959_ (.A1(_3311_),
    .A2(_3248_),
    .B(_3312_),
    .C(_0904_),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7960_ (.A1(_2050_),
    .A2(_3162_),
    .B(_3159_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7961_ (.A1(_2156_),
    .A2(_2976_),
    .B(_3314_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7962_ (.A1(_1561_),
    .A2(_1361_),
    .B1(_3313_),
    .B2(_3315_),
    .C(_1684_),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7963_ (.A1(_1644_),
    .A2(_3316_),
    .B(_3274_),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7964_ (.A1(_1741_),
    .A2(_1643_),
    .B(_3317_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7965_ (.A1(_0878_),
    .A2(_3198_),
    .B1(_1623_),
    .B2(_1624_),
    .C(_3318_),
    .ZN(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7966_ (.A1(_3310_),
    .A2(_3319_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7967_ (.I(_2581_),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7968_ (.A1(_1059_),
    .A2(_3197_),
    .B(_3321_),
    .ZN(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7969_ (.A1(_3203_),
    .A2(_3320_),
    .B(_3322_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7970_ (.A1(_1112_),
    .A2(_1183_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7971_ (.I(_3323_),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7972_ (.I(_3324_),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7973_ (.I(_3323_),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7974_ (.I(_3326_),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7975_ (.A1(\as2650.stack[7][8] ),
    .A2(_3327_),
    .ZN(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7976_ (.A1(_1478_),
    .A2(_3325_),
    .B(_3328_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7977_ (.I(_3326_),
    .Z(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7978_ (.A1(\as2650.stack[7][9] ),
    .A2(_3329_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7979_ (.A1(_1487_),
    .A2(_3325_),
    .B(_3330_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7980_ (.A1(\as2650.stack[7][10] ),
    .A2(_3329_),
    .ZN(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7981_ (.A1(_1490_),
    .A2(_3325_),
    .B(_3331_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7982_ (.A1(\as2650.stack[7][11] ),
    .A2(_3329_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7983_ (.A1(_1492_),
    .A2(_3325_),
    .B(_3332_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7984_ (.I(_3324_),
    .Z(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7985_ (.A1(\as2650.stack[7][12] ),
    .A2(_3329_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7986_ (.A1(_1494_),
    .A2(_3333_),
    .B(_3334_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7987_ (.I(_3326_),
    .Z(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7988_ (.A1(\as2650.stack[7][13] ),
    .A2(_3335_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7989_ (.A1(_1497_),
    .A2(_3333_),
    .B(_3336_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7990_ (.A1(\as2650.stack[7][14] ),
    .A2(_3335_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7991_ (.A1(_1500_),
    .A2(_3333_),
    .B(_3337_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7992_ (.I(_1185_),
    .Z(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7993_ (.I(_3338_),
    .Z(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7994_ (.A1(\as2650.stack[6][0] ),
    .A2(_1231_),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7995_ (.A1(_2116_),
    .A2(_3339_),
    .B(_3340_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7996_ (.A1(\as2650.stack[6][1] ),
    .A2(_1231_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7997_ (.A1(_2123_),
    .A2(_3339_),
    .B(_3341_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7998_ (.I(_1185_),
    .Z(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7999_ (.A1(\as2650.stack[6][2] ),
    .A2(_3342_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8000_ (.A1(_2126_),
    .A2(_3339_),
    .B(_3343_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8001_ (.A1(\as2650.stack[6][3] ),
    .A2(_3342_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8002_ (.A1(_2128_),
    .A2(_3339_),
    .B(_3344_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8003_ (.I(_3338_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8004_ (.A1(\as2650.stack[6][4] ),
    .A2(_3342_),
    .ZN(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8005_ (.A1(_2130_),
    .A2(_3345_),
    .B(_3346_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8006_ (.A1(\as2650.stack[6][5] ),
    .A2(_3342_),
    .ZN(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8007_ (.A1(_2133_),
    .A2(_3345_),
    .B(_3347_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8008_ (.A1(\as2650.stack[6][6] ),
    .A2(_3338_),
    .ZN(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8009_ (.A1(_2136_),
    .A2(_3345_),
    .B(_3348_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8010_ (.A1(\as2650.stack[6][7] ),
    .A2(_3338_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8011_ (.A1(_2138_),
    .A2(_3345_),
    .B(_3349_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8012_ (.I(_1122_),
    .Z(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8013_ (.A1(\as2650.stack[5][8] ),
    .A2(_1165_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8014_ (.A1(_3350_),
    .A2(_1193_),
    .B(_3351_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8015_ (.I(_1113_),
    .Z(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8016_ (.A1(\as2650.stack[5][9] ),
    .A2(_3352_),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8017_ (.A1(_3350_),
    .A2(_1201_),
    .B(_3353_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8018_ (.A1(\as2650.stack[5][10] ),
    .A2(_3352_),
    .ZN(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8019_ (.A1(_3350_),
    .A2(_1208_),
    .B(_3354_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8020_ (.A1(\as2650.stack[5][11] ),
    .A2(_3352_),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8021_ (.A1(_3350_),
    .A2(_1217_),
    .B(_3355_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8022_ (.A1(\as2650.stack[5][12] ),
    .A2(_3352_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8023_ (.A1(_1123_),
    .A2(_1224_),
    .B(_3356_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8024_ (.A1(\as2650.stack[5][13] ),
    .A2(_1114_),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8025_ (.A1(_1123_),
    .A2(_1230_),
    .B(_3357_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8026_ (.A1(\as2650.stack[5][14] ),
    .A2(_1114_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8027_ (.A1(_1123_),
    .A2(_1237_),
    .B(_3358_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8028_ (.I(_2120_),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8029_ (.A1(\as2650.stack[4][8] ),
    .A2(_2134_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8030_ (.A1(_1478_),
    .A2(_3359_),
    .B(_3360_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8031_ (.I(_2117_),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8032_ (.A1(\as2650.stack[4][9] ),
    .A2(_3361_),
    .ZN(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8033_ (.A1(_1487_),
    .A2(_3359_),
    .B(_3362_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8034_ (.A1(\as2650.stack[4][10] ),
    .A2(_3361_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8035_ (.A1(_1490_),
    .A2(_3359_),
    .B(_3363_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8036_ (.A1(\as2650.stack[4][11] ),
    .A2(_3361_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8037_ (.A1(_1492_),
    .A2(_3359_),
    .B(_3364_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8038_ (.A1(\as2650.stack[4][12] ),
    .A2(_3361_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8039_ (.A1(_1494_),
    .A2(_2121_),
    .B(_3365_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8040_ (.A1(\as2650.stack[4][13] ),
    .A2(_2118_),
    .ZN(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8041_ (.A1(_1497_),
    .A2(_2121_),
    .B(_3366_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8042_ (.A1(\as2650.stack[4][14] ),
    .A2(_2118_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8043_ (.A1(_1500_),
    .A2(_2121_),
    .B(_3367_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8044_ (.A1(\as2650.stack[7][0] ),
    .A2(_3335_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8045_ (.A1(_2116_),
    .A2(_3333_),
    .B(_3368_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8046_ (.I(_3326_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8047_ (.A1(\as2650.stack[7][1] ),
    .A2(_3335_),
    .ZN(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8048_ (.A1(_2123_),
    .A2(_3369_),
    .B(_3370_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8049_ (.I(_3323_),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8050_ (.A1(\as2650.stack[7][2] ),
    .A2(_3371_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8051_ (.A1(_2126_),
    .A2(_3369_),
    .B(_3372_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8052_ (.A1(\as2650.stack[7][3] ),
    .A2(_3371_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8053_ (.A1(_2128_),
    .A2(_3369_),
    .B(_3373_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8054_ (.A1(\as2650.stack[7][4] ),
    .A2(_3371_),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8055_ (.A1(_2130_),
    .A2(_3369_),
    .B(_3374_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8056_ (.A1(\as2650.stack[7][5] ),
    .A2(_3371_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8057_ (.A1(_2133_),
    .A2(_3327_),
    .B(_3375_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8058_ (.A1(\as2650.stack[7][6] ),
    .A2(_3324_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8059_ (.A1(_2136_),
    .A2(_3327_),
    .B(_3376_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8060_ (.A1(\as2650.stack[7][7] ),
    .A2(_3324_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8061_ (.A1(_2138_),
    .A2(_3327_),
    .B(_3377_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8062_ (.A1(_0851_),
    .A2(_1597_),
    .A3(_1616_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8063_ (.A1(_1614_),
    .A2(_3378_),
    .ZN(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8064_ (.A1(_2653_),
    .A2(_2312_),
    .B(_2317_),
    .C(_3379_),
    .ZN(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8065_ (.A1(_2241_),
    .A2(_2322_),
    .A3(_2341_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8066_ (.A1(_2159_),
    .A2(_2592_),
    .A3(_3380_),
    .A4(_3381_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8067_ (.A1(_2223_),
    .A2(_2237_),
    .B(_2312_),
    .ZN(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8068_ (.A1(_1241_),
    .A2(_2818_),
    .A3(_1249_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8069_ (.A1(_3383_),
    .A2(_3384_),
    .B(_1429_),
    .C(_2229_),
    .ZN(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8070_ (.A1(_2339_),
    .A2(_2589_),
    .A3(_3382_),
    .A4(_3385_),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8071_ (.A1(_2311_),
    .A2(_3386_),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8072_ (.I(_3387_),
    .Z(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8073_ (.I(_3388_),
    .Z(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8074_ (.I(_3389_),
    .Z(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8075_ (.I(_1314_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8076_ (.A1(_3191_),
    .A2(_4062_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8077_ (.A1(_1530_),
    .A2(_3392_),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8078_ (.A1(_3978_),
    .A2(_4131_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8079_ (.A1(_2632_),
    .A2(_3394_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8080_ (.I(_1322_),
    .Z(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8081_ (.I(_3396_),
    .Z(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8082_ (.I(_3397_),
    .Z(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8083_ (.A1(_2564_),
    .A2(_3393_),
    .B1(_3395_),
    .B2(_3398_),
    .ZN(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8084_ (.I(net28),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8085_ (.A1(_3911_),
    .A2(_1294_),
    .Z(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8086_ (.I(_3401_),
    .Z(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8087_ (.A1(_3400_),
    .A2(_3402_),
    .B1(_2484_),
    .B2(_2612_),
    .C(_1318_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8088_ (.A1(_3391_),
    .A2(_3399_),
    .B(_3403_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8089_ (.A1(_1395_),
    .A2(_2945_),
    .B(_2301_),
    .ZN(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8090_ (.I(_3405_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8091_ (.A1(_2678_),
    .A2(_2337_),
    .ZN(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8092_ (.I(_3407_),
    .Z(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8093_ (.A1(_2632_),
    .A2(_2734_),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8094_ (.A1(_3400_),
    .A2(_2829_),
    .B(_3409_),
    .ZN(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8095_ (.A1(_2505_),
    .A2(_2612_),
    .B1(_3408_),
    .B2(_3410_),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8096_ (.I(_2719_),
    .Z(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8097_ (.A1(_1119_),
    .A2(_3406_),
    .B1(_3411_),
    .B2(_3412_),
    .ZN(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8098_ (.A1(_1571_),
    .A2(_3413_),
    .ZN(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8099_ (.A1(_3404_),
    .A2(_3414_),
    .ZN(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8100_ (.A1(_3221_),
    .A2(_2299_),
    .ZN(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8101_ (.A1(_2353_),
    .A2(_3415_),
    .B1(_3416_),
    .B2(_2609_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8102_ (.I(_3388_),
    .Z(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8103_ (.A1(_3400_),
    .A2(_3418_),
    .B(_3321_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8104_ (.A1(_3390_),
    .A2(_3417_),
    .B(_3419_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8105_ (.A1(_1622_),
    .A2(_2287_),
    .ZN(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8106_ (.I(_3420_),
    .Z(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8107_ (.I(_3421_),
    .Z(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8108_ (.I(_1295_),
    .Z(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8109_ (.A1(net52),
    .A2(_3400_),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8110_ (.I(_1315_),
    .Z(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8111_ (.A1(_2486_),
    .A2(_3921_),
    .ZN(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8112_ (.I(_3426_),
    .Z(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _8113_ (.A1(_4068_),
    .A2(_4061_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _8114_ (.A1(_2250_),
    .A2(_4238_),
    .A3(_4241_),
    .Z(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8115_ (.A1(_3428_),
    .A2(_3429_),
    .Z(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8116_ (.A1(_1321_),
    .A2(_3191_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8117_ (.I(_3431_),
    .Z(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8118_ (.I(_3189_),
    .Z(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8119_ (.A1(_4068_),
    .A2(_4130_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8120_ (.A1(_2251_),
    .A2(_4236_),
    .A3(_3434_),
    .Z(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8121_ (.I(_4123_),
    .Z(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8122_ (.A1(_4272_),
    .A2(_3436_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8123_ (.A1(_3433_),
    .A2(_3435_),
    .B(_3437_),
    .C(_3397_),
    .ZN(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8124_ (.A1(_4272_),
    .A2(_3427_),
    .B1(_3430_),
    .B2(_3432_),
    .C(_3438_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8125_ (.A1(_3425_),
    .A2(_3439_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8126_ (.I(_2407_),
    .Z(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8127_ (.A1(_3423_),
    .A2(_3424_),
    .B(_3440_),
    .C(_3441_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8128_ (.I(_2483_),
    .Z(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8129_ (.A1(_1116_),
    .A2(_4068_),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8130_ (.A1(_3444_),
    .A2(_2670_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8131_ (.A1(_3443_),
    .A2(_3445_),
    .B(_3281_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8132_ (.A1(_2734_),
    .A2(_3424_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8133_ (.A1(_2680_),
    .A2(_3447_),
    .Z(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8134_ (.A1(_3132_),
    .A2(_2671_),
    .B1(_3408_),
    .B2(_3448_),
    .ZN(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8135_ (.A1(_2669_),
    .A2(_3406_),
    .B1(_3449_),
    .B2(_3412_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8136_ (.A1(_3442_),
    .A2(_3446_),
    .B1(_3450_),
    .B2(_1571_),
    .ZN(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8137_ (.I(_2287_),
    .Z(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8138_ (.I(_3452_),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8139_ (.A1(_2669_),
    .A2(_3422_),
    .B1(_3451_),
    .B2(_3453_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8140_ (.A1(net52),
    .A2(_3418_),
    .B(_3321_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8141_ (.A1(_3390_),
    .A2(_3454_),
    .B(_3455_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8142_ (.I(_3978_),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8143_ (.A1(_4232_),
    .A2(_4235_),
    .B(_4269_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8144_ (.A1(_4269_),
    .A2(_4232_),
    .A3(_4235_),
    .ZN(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8145_ (.A1(_3434_),
    .A2(_3457_),
    .B(_3458_),
    .ZN(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8146_ (.A1(_0389_),
    .A2(_0392_),
    .B(_1663_),
    .ZN(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8147_ (.A1(_0353_),
    .A2(_0393_),
    .ZN(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8148_ (.A1(_3460_),
    .A2(_3461_),
    .ZN(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8149_ (.A1(_3459_),
    .A2(_3462_),
    .B(_3433_),
    .ZN(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8150_ (.A1(_3459_),
    .A2(_3462_),
    .B(_3463_),
    .ZN(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8151_ (.A1(_1532_),
    .A2(_3456_),
    .B(_3398_),
    .C(_3464_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _8152_ (.A1(_2250_),
    .A2(_4242_),
    .A3(_4243_),
    .B1(_3428_),
    .B2(_3429_),
    .ZN(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8153_ (.A1(_2255_),
    .A2(_0386_),
    .A3(_3466_),
    .Z(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8154_ (.A1(_1532_),
    .A2(_3192_),
    .B1(_3467_),
    .B2(_3922_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8155_ (.A1(_3465_),
    .A2(_3468_),
    .ZN(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8156_ (.A1(_2404_),
    .A2(_3469_),
    .ZN(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8157_ (.A1(net52),
    .A2(net28),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8158_ (.A1(net30),
    .A2(_3471_),
    .ZN(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8159_ (.A1(_3444_),
    .A2(_2713_),
    .B(_2714_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8160_ (.A1(_2717_),
    .A2(_3473_),
    .Z(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8161_ (.A1(_3402_),
    .A2(_3472_),
    .B1(_3474_),
    .B2(_3443_),
    .ZN(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8162_ (.A1(_3470_),
    .A2(_3475_),
    .B(_3155_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8163_ (.A1(_2876_),
    .A2(_3472_),
    .B(_2725_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8164_ (.A1(_2505_),
    .A2(_2718_),
    .B1(_3408_),
    .B2(_3477_),
    .ZN(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8165_ (.A1(_1137_),
    .A2(_3406_),
    .B1(_3478_),
    .B2(_3412_),
    .ZN(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8166_ (.I(_3387_),
    .Z(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8167_ (.A1(_1139_),
    .A2(_3421_),
    .B1(_3479_),
    .B2(_2661_),
    .C(_3480_),
    .ZN(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8168_ (.A1(_2353_),
    .A2(_3476_),
    .B(_3481_),
    .ZN(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8169_ (.I(_3480_),
    .Z(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8170_ (.A1(net30),
    .A2(_3483_),
    .B(_3224_),
    .ZN(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8171_ (.A1(_3482_),
    .A2(_3484_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8172_ (.I(_3480_),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8173_ (.I(_3420_),
    .Z(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8174_ (.A1(net30),
    .A2(net29),
    .A3(net28),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8175_ (.A1(net31),
    .A2(_3487_),
    .Z(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8176_ (.A1(_3401_),
    .A2(_3488_),
    .B(_2484_),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8177_ (.A1(_1954_),
    .A2(_0385_),
    .ZN(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8178_ (.A1(_1663_),
    .A2(_0385_),
    .ZN(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8179_ (.A1(_3466_),
    .A2(_3490_),
    .B(_3491_),
    .ZN(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8180_ (.A1(_0426_),
    .A2(_0454_),
    .A3(_3492_),
    .ZN(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8181_ (.A1(_1663_),
    .A2(_0389_),
    .A3(_0392_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8182_ (.A1(_3459_),
    .A2(_3460_),
    .B(_3494_),
    .ZN(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8183_ (.A1(_0425_),
    .A2(_0459_),
    .A3(_3495_),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8184_ (.A1(_0427_),
    .A2(_3436_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8185_ (.A1(_3433_),
    .A2(_3496_),
    .B(_3497_),
    .C(_3396_),
    .ZN(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8186_ (.A1(_1533_),
    .A2(_3427_),
    .B1(_3493_),
    .B2(_3432_),
    .C(_3498_),
    .ZN(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8187_ (.A1(_1315_),
    .A2(_3499_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8188_ (.A1(_2717_),
    .A2(_3473_),
    .ZN(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8189_ (.A1(_2762_),
    .A2(_3501_),
    .ZN(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8190_ (.A1(_2761_),
    .A2(_3502_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8191_ (.A1(_3489_),
    .A2(_3500_),
    .B1(_3503_),
    .B2(_3443_),
    .ZN(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8192_ (.A1(_1396_),
    .A2(_2945_),
    .ZN(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8193_ (.I(_3407_),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8194_ (.A1(_2293_),
    .A2(_3488_),
    .B(_2769_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8195_ (.A1(_2323_),
    .A2(_3506_),
    .A3(_3507_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8196_ (.A1(_2946_),
    .A2(_2765_),
    .B1(_3505_),
    .B2(_1145_),
    .C(_3508_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8197_ (.A1(_1720_),
    .A2(_3509_),
    .ZN(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8198_ (.A1(_1145_),
    .A2(_3274_),
    .B1(_3226_),
    .B2(_3504_),
    .C(_3510_),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8199_ (.A1(_2757_),
    .A2(_3486_),
    .B1(_3511_),
    .B2(_3452_),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8200_ (.A1(net31),
    .A2(_3389_),
    .ZN(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8201_ (.A1(_3485_),
    .A2(_3512_),
    .B(_3513_),
    .C(_3135_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8202_ (.A1(_2824_),
    .A2(_0459_),
    .ZN(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _8203_ (.A1(_2824_),
    .A2(_0459_),
    .B1(_3459_),
    .B2(_3460_),
    .C(_3494_),
    .ZN(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8204_ (.A1(_3514_),
    .A2(_3515_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8205_ (.A1(_1660_),
    .A2(_0556_),
    .A3(_3516_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8206_ (.A1(_3456_),
    .A2(_3517_),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8207_ (.A1(_0561_),
    .A2(_3456_),
    .B(_3397_),
    .C(_3518_),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8208_ (.A1(_0424_),
    .A2(_0453_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _8209_ (.A1(_0424_),
    .A2(_0453_),
    .B1(_3466_),
    .B2(_3490_),
    .C(_3491_),
    .ZN(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8210_ (.A1(_3520_),
    .A2(_3521_),
    .ZN(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8211_ (.A1(_2031_),
    .A2(_0594_),
    .A3(_3522_),
    .Z(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8212_ (.A1(_0561_),
    .A2(_3192_),
    .B1(_3523_),
    .B2(_3922_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8213_ (.A1(_3519_),
    .A2(_3524_),
    .B(_1314_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8214_ (.A1(_2757_),
    .A2(_2824_),
    .Z(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8215_ (.A1(_2760_),
    .A2(_3502_),
    .Z(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8216_ (.A1(_3526_),
    .A2(_2808_),
    .A3(_3527_),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8217_ (.A1(_3526_),
    .A2(_3527_),
    .B(_2808_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8218_ (.I(net31),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8219_ (.A1(_3530_),
    .A2(_3487_),
    .ZN(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8220_ (.A1(net32),
    .A2(_3531_),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8221_ (.A1(_2408_),
    .A2(_3528_),
    .A3(_3529_),
    .B1(_3532_),
    .B2(_3423_),
    .ZN(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8222_ (.A1(_3525_),
    .A2(_3533_),
    .B(_2300_),
    .C(_3226_),
    .ZN(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8223_ (.A1(_1269_),
    .A2(_3532_),
    .B(_2819_),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8224_ (.A1(_2777_),
    .A2(_2811_),
    .B1(_3506_),
    .B2(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8225_ (.A1(_1152_),
    .A2(_3405_),
    .B1(_3536_),
    .B2(_2720_),
    .C(_2660_),
    .ZN(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8226_ (.A1(_2857_),
    .A2(_3416_),
    .B(_3537_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8227_ (.A1(_3480_),
    .A2(_3534_),
    .A3(_3538_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8228_ (.A1(net32),
    .A2(_3483_),
    .B(_3539_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8229_ (.A1(_3242_),
    .A2(_3540_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8230_ (.I(_2408_),
    .Z(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8231_ (.A1(_3526_),
    .A2(_2808_),
    .A3(_3527_),
    .ZN(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8232_ (.A1(_2906_),
    .A2(_3542_),
    .ZN(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8233_ (.A1(_2856_),
    .A2(_3543_),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8234_ (.A1(net32),
    .A2(_3531_),
    .Z(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8235_ (.A1(net51),
    .A2(_3545_),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8236_ (.A1(_1674_),
    .A2(_0593_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8237_ (.A1(_0560_),
    .A2(_0593_),
    .ZN(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _8238_ (.A1(_3520_),
    .A2(_3547_),
    .A3(_3521_),
    .B(_3548_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8239_ (.A1(_0657_),
    .A2(_0682_),
    .A3(_3549_),
    .Z(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8240_ (.A1(_0657_),
    .A2(_0654_),
    .Z(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8241_ (.A1(_1674_),
    .A2(_0555_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8242_ (.A1(_1674_),
    .A2(_0555_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _8243_ (.A1(_3514_),
    .A2(_3552_),
    .A3(_3515_),
    .B(_3553_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8244_ (.A1(_3551_),
    .A2(_3554_),
    .B(_3189_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8245_ (.A1(_3551_),
    .A2(_3554_),
    .B(_3555_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8246_ (.A1(_2063_),
    .A2(_3456_),
    .B(_3397_),
    .C(_3556_),
    .ZN(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8247_ (.A1(_0658_),
    .A2(_3427_),
    .B1(_3550_),
    .B2(_3432_),
    .C(_3557_),
    .ZN(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8248_ (.A1(_3402_),
    .A2(_3546_),
    .B1(_3558_),
    .B2(_3425_),
    .ZN(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8249_ (.A1(_3441_),
    .A2(_3559_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8250_ (.A1(_3541_),
    .A2(_3544_),
    .B(_3560_),
    .C(_3296_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8251_ (.I(_2330_),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8252_ (.I(_2391_),
    .Z(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8253_ (.A1(_3563_),
    .A2(_3546_),
    .B(_2866_),
    .ZN(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8254_ (.A1(_2898_),
    .A2(_2297_),
    .B1(_3562_),
    .B2(_3564_),
    .ZN(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8255_ (.A1(_2992_),
    .A2(_2666_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8256_ (.I(_3566_),
    .Z(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8257_ (.A1(_2898_),
    .A2(_3567_),
    .B(_2664_),
    .ZN(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8258_ (.A1(_2863_),
    .A2(_2861_),
    .B1(_3565_),
    .B2(_1736_),
    .C(_3568_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8259_ (.A1(_2898_),
    .A2(_3422_),
    .B1(_3561_),
    .B2(_3453_),
    .C(_3569_),
    .ZN(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8260_ (.A1(net51),
    .A2(_3418_),
    .B(_3321_),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8261_ (.A1(_3390_),
    .A2(_3570_),
    .B(_3571_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8262_ (.A1(net51),
    .A2(_3545_),
    .ZN(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8263_ (.A1(net34),
    .A2(_3572_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8264_ (.A1(_0730_),
    .A2(_0725_),
    .Z(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8265_ (.I(_0656_),
    .Z(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8266_ (.A1(_3575_),
    .A2(_0681_),
    .Z(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8267_ (.A1(_3575_),
    .A2(_0681_),
    .Z(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8268_ (.A1(_3576_),
    .A2(_3549_),
    .B(_3577_),
    .ZN(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8269_ (.A1(_3574_),
    .A2(_3578_),
    .Z(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8270_ (.A1(_3575_),
    .A2(_0653_),
    .Z(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8271_ (.A1(_3575_),
    .A2(_0653_),
    .Z(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _8272_ (.A1(_3580_),
    .A2(_3554_),
    .B(_3581_),
    .ZN(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8273_ (.A1(_2084_),
    .A2(_0722_),
    .A3(_3582_),
    .Z(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8274_ (.A1(_1539_),
    .A2(_3436_),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8275_ (.A1(_3433_),
    .A2(_3583_),
    .B(_3584_),
    .C(_3396_),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8276_ (.A1(_1541_),
    .A2(_3427_),
    .B1(_3579_),
    .B2(_3432_),
    .C(_3585_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8277_ (.A1(_3425_),
    .A2(_3586_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8278_ (.I(_2407_),
    .Z(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8279_ (.A1(_3423_),
    .A2(_3573_),
    .B(_3587_),
    .C(_3588_),
    .ZN(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _8280_ (.A1(_2855_),
    .A2(_2907_),
    .B1(_3528_),
    .B2(_2856_),
    .ZN(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8281_ (.A1(_2904_),
    .A2(_3590_),
    .Z(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8282_ (.A1(_3443_),
    .A2(_3591_),
    .B(_3281_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8283_ (.A1(_2228_),
    .A2(_3573_),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8284_ (.A1(_2920_),
    .A2(_3593_),
    .Z(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8285_ (.A1(_2777_),
    .A2(_2910_),
    .B1(_3506_),
    .B2(_3594_),
    .ZN(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8286_ (.A1(_1168_),
    .A2(_3405_),
    .B1(_3595_),
    .B2(_2720_),
    .ZN(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8287_ (.A1(_3589_),
    .A2(_3592_),
    .B1(_3596_),
    .B2(_2279_),
    .ZN(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8288_ (.A1(_1168_),
    .A2(_3486_),
    .B1(_3597_),
    .B2(_3452_),
    .ZN(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8289_ (.A1(net34),
    .A2(_3389_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8290_ (.A1(_3483_),
    .A2(_3598_),
    .B(_3599_),
    .C(_3135_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8291_ (.A1(_2904_),
    .A2(_3590_),
    .B(_2948_),
    .ZN(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8292_ (.A1(_2947_),
    .A2(_3600_),
    .ZN(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8293_ (.A1(_1538_),
    .A2(_0726_),
    .ZN(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8294_ (.A1(_3574_),
    .A2(_3578_),
    .B(_3602_),
    .ZN(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8295_ (.A1(_1647_),
    .A2(_0886_),
    .A3(_3603_),
    .Z(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8296_ (.A1(_1538_),
    .A2(_0721_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8297_ (.A1(_1538_),
    .A2(_0721_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8298_ (.A1(_3605_),
    .A2(_3582_),
    .B(_3606_),
    .ZN(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8299_ (.A1(_0875_),
    .A2(_2104_),
    .A3(_3607_),
    .Z(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8300_ (.A1(_0876_),
    .A2(_3189_),
    .ZN(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8301_ (.A1(_3436_),
    .A2(_3608_),
    .B(_3609_),
    .C(_3396_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8302_ (.A1(_1543_),
    .A2(_3426_),
    .B1(_3604_),
    .B2(_3431_),
    .C(_3610_),
    .ZN(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8303_ (.A1(net34),
    .A2(net51),
    .A3(_3545_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8304_ (.A1(net35),
    .A2(_3612_),
    .Z(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8305_ (.A1(_1315_),
    .A2(_3611_),
    .B1(_3613_),
    .B2(_3401_),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8306_ (.A1(_3441_),
    .A2(_3614_),
    .ZN(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8307_ (.A1(_3541_),
    .A2(_3601_),
    .B(_3615_),
    .C(_1524_),
    .ZN(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8308_ (.A1(_1543_),
    .A2(_2460_),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8309_ (.A1(_3563_),
    .A2(_3613_),
    .B(_3617_),
    .ZN(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8310_ (.A1(_2994_),
    .A2(_2297_),
    .B1(_3562_),
    .B2(_3618_),
    .ZN(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8311_ (.A1(_2994_),
    .A2(_3566_),
    .B(_2660_),
    .ZN(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8312_ (.A1(_2389_),
    .A2(_3619_),
    .B(_3620_),
    .C(_2952_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8313_ (.A1(_2994_),
    .A2(_3421_),
    .B1(_3616_),
    .B2(_3452_),
    .C(_3621_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8314_ (.A1(net35),
    .A2(_3389_),
    .ZN(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8315_ (.I(_2414_),
    .Z(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8316_ (.A1(_3483_),
    .A2(_3622_),
    .B(_3623_),
    .C(_3624_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8317_ (.A1(_0875_),
    .A2(_0885_),
    .ZN(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _8318_ (.A1(_3574_),
    .A2(_3578_),
    .B(_3625_),
    .C(_3602_),
    .ZN(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8319_ (.A1(_0875_),
    .A2(_0885_),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8320_ (.A1(_3921_),
    .A2(_3627_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8321_ (.A1(_3626_),
    .A2(_3628_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8322_ (.A1(_2247_),
    .A2(_3629_),
    .Z(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _8323_ (.A1(_1300_),
    .A2(_2104_),
    .B1(_3605_),
    .B2(_3582_),
    .C(_3606_),
    .ZN(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8324_ (.A1(_1300_),
    .A2(_2104_),
    .B(_4123_),
    .ZN(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8325_ (.A1(_3631_),
    .A2(_3632_),
    .ZN(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8326_ (.A1(_2247_),
    .A2(_3633_),
    .Z(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8327_ (.A1(_2564_),
    .A2(_3630_),
    .B1(_3634_),
    .B2(_3398_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8328_ (.I(net36),
    .Z(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8329_ (.I(net35),
    .ZN(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8330_ (.A1(_3637_),
    .A2(_3612_),
    .ZN(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8331_ (.A1(_3636_),
    .A2(_3638_),
    .Z(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8332_ (.A1(_3423_),
    .A2(_3639_),
    .Z(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8333_ (.A1(_3391_),
    .A2(_3635_),
    .B(_3640_),
    .C(_3441_),
    .ZN(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8334_ (.A1(_2984_),
    .A2(_3590_),
    .B(_2986_),
    .ZN(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8335_ (.A1(_2983_),
    .A2(_3642_),
    .Z(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8336_ (.A1(_3588_),
    .A2(_3643_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8337_ (.A1(_2983_),
    .A2(_3642_),
    .B(_3644_),
    .ZN(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8338_ (.A1(_2300_),
    .A2(_1525_),
    .A3(_3641_),
    .A4(_3645_),
    .ZN(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8339_ (.A1(_2470_),
    .A2(_3505_),
    .ZN(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8340_ (.A1(_2471_),
    .A2(_3639_),
    .ZN(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8341_ (.A1(_2247_),
    .A2(_2460_),
    .B(_3506_),
    .ZN(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8342_ (.A1(_2529_),
    .A2(_2989_),
    .B1(_3648_),
    .B2(_3649_),
    .ZN(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8343_ (.A1(_1190_),
    .A2(_3647_),
    .B1(_3650_),
    .B2(_3567_),
    .ZN(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8344_ (.A1(_2656_),
    .A2(_3651_),
    .ZN(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8345_ (.A1(_1190_),
    .A2(_3422_),
    .B(_3646_),
    .C(_3652_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8346_ (.I(_3388_),
    .Z(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8347_ (.I(_3903_),
    .Z(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8348_ (.A1(_3636_),
    .A2(_3654_),
    .B(_3655_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8349_ (.A1(_3390_),
    .A2(_3653_),
    .B(_3656_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8350_ (.A1(_1189_),
    .A2(_1540_),
    .B(_3643_),
    .ZN(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8351_ (.A1(_3018_),
    .A2(_3657_),
    .Z(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8352_ (.A1(_3001_),
    .A2(_3631_),
    .A3(_3632_),
    .ZN(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8353_ (.A1(_2252_),
    .A2(_3659_),
    .Z(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8354_ (.A1(_3001_),
    .A2(_3626_),
    .A3(_3628_),
    .ZN(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8355_ (.A1(_2252_),
    .A2(_3661_),
    .Z(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8356_ (.A1(_3398_),
    .A2(_3660_),
    .B1(_3662_),
    .B2(_2569_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8357_ (.A1(_3636_),
    .A2(_3638_),
    .ZN(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8358_ (.A1(net50),
    .A2(_3664_),
    .Z(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8359_ (.A1(_3402_),
    .A2(_3665_),
    .ZN(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8360_ (.A1(_3391_),
    .A2(_3663_),
    .B(_3666_),
    .C(_3588_),
    .ZN(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8361_ (.A1(_3541_),
    .A2(_3658_),
    .B(_3667_),
    .C(_3296_),
    .ZN(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8362_ (.A1(_2481_),
    .A2(_3665_),
    .B(_3032_),
    .ZN(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8363_ (.A1(_3028_),
    .A2(_2283_),
    .B1(_3562_),
    .B2(_3669_),
    .ZN(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8364_ (.A1(_3028_),
    .A2(_3567_),
    .B(_2664_),
    .ZN(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8365_ (.A1(_1736_),
    .A2(_3670_),
    .B(_3671_),
    .C(_3023_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8366_ (.A1(_3028_),
    .A2(_3486_),
    .B1(_3668_),
    .B2(_3453_),
    .C(_3672_),
    .ZN(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8367_ (.A1(net50),
    .A2(_3654_),
    .B(_3655_),
    .ZN(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8368_ (.A1(_3485_),
    .A2(_3673_),
    .B(_3674_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8369_ (.A1(net50),
    .A2(_3636_),
    .A3(_3638_),
    .ZN(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8370_ (.A1(net38),
    .A2(_3675_),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8371_ (.A1(_2876_),
    .A2(_3676_),
    .B(_3060_),
    .ZN(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8372_ (.A1(_3132_),
    .A2(_3050_),
    .B1(_3408_),
    .B2(_3677_),
    .ZN(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8373_ (.A1(_3042_),
    .A2(_3406_),
    .B1(_3678_),
    .B2(_3412_),
    .C(_1688_),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8374_ (.A1(_3018_),
    .A2(_3643_),
    .Z(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8375_ (.A1(_3048_),
    .A2(_3680_),
    .ZN(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8376_ (.A1(_3044_),
    .A2(_3681_),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8377_ (.A1(_1240_),
    .A2(_1295_),
    .Z(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8378_ (.A1(_3631_),
    .A2(_3632_),
    .B(_1321_),
    .ZN(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8379_ (.A1(_2630_),
    .A2(_2252_),
    .B(_1297_),
    .ZN(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8380_ (.A1(_3626_),
    .A2(_3628_),
    .B(_2216_),
    .ZN(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8381_ (.A1(_3683_),
    .A2(_3684_),
    .B(_3685_),
    .C(_3686_),
    .ZN(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _8382_ (.A1(_1296_),
    .A2(_3075_),
    .A3(_3686_),
    .A4(_3684_),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8383_ (.A1(_2256_),
    .A2(_3687_),
    .B(_3688_),
    .ZN(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8384_ (.A1(_1295_),
    .A2(_3676_),
    .B(_2407_),
    .ZN(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8385_ (.A1(_2404_),
    .A2(_3689_),
    .B(_3690_),
    .ZN(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8386_ (.A1(_2544_),
    .A2(_3682_),
    .B(_3691_),
    .C(_3281_),
    .ZN(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8387_ (.A1(_3679_),
    .A2(_3692_),
    .B(_2400_),
    .ZN(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8388_ (.A1(_3042_),
    .A2(_3422_),
    .B(_3693_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8389_ (.A1(net38),
    .A2(_3654_),
    .B(_3655_),
    .ZN(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8390_ (.A1(_3485_),
    .A2(_3694_),
    .B(_3695_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8391_ (.I(_3088_),
    .Z(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8392_ (.A1(_3044_),
    .A2(_3681_),
    .B(_3081_),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8393_ (.A1(_3080_),
    .A2(_3697_),
    .Z(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8394_ (.A1(_3683_),
    .A2(_3075_),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _8395_ (.A1(_3683_),
    .A2(_3684_),
    .B(_3699_),
    .C(_3686_),
    .ZN(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8396_ (.I(_2259_),
    .ZN(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8397_ (.I0(_3688_),
    .I1(_3700_),
    .S(_3701_),
    .Z(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8398_ (.A1(net38),
    .A2(net50),
    .A3(net36),
    .A4(_3638_),
    .ZN(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8399_ (.A1(net39),
    .A2(_3703_),
    .Z(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8400_ (.A1(_3401_),
    .A2(_3704_),
    .ZN(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8401_ (.A1(_1314_),
    .A2(_3702_),
    .B(_3705_),
    .C(_3588_),
    .ZN(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8402_ (.A1(_3541_),
    .A2(_3698_),
    .B(_3706_),
    .C(_3296_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8403_ (.A1(_3563_),
    .A2(_3704_),
    .B(_3084_),
    .ZN(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8404_ (.A1(_3696_),
    .A2(_2297_),
    .B1(_3562_),
    .B2(_3708_),
    .ZN(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8405_ (.A1(_3696_),
    .A2(_3567_),
    .B(_2664_),
    .ZN(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8406_ (.A1(_2863_),
    .A2(_3083_),
    .B1(_3709_),
    .B2(_2389_),
    .C(_3710_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8407_ (.A1(_3696_),
    .A2(_3486_),
    .B1(_3707_),
    .B2(_3453_),
    .C(_3711_),
    .ZN(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8408_ (.A1(net39),
    .A2(_3654_),
    .B(_3655_),
    .ZN(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8409_ (.A1(_3485_),
    .A2(_3712_),
    .B(_3713_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8410_ (.A1(_3696_),
    .A2(_1540_),
    .B1(_3101_),
    .B2(_3680_),
    .C(_3102_),
    .ZN(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8411_ (.A1(_3104_),
    .A2(_3714_),
    .Z(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8412_ (.I(net39),
    .ZN(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8413_ (.A1(_3716_),
    .A2(_3703_),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8414_ (.A1(net40),
    .A2(_3717_),
    .ZN(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8415_ (.A1(_3701_),
    .A2(_3688_),
    .B(_2261_),
    .ZN(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8416_ (.A1(_2259_),
    .A2(_1297_),
    .B(_3700_),
    .C(_2817_),
    .ZN(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8417_ (.A1(_1297_),
    .A2(_3718_),
    .B1(_3719_),
    .B2(_3720_),
    .ZN(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8418_ (.A1(_2558_),
    .A2(_3718_),
    .ZN(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8419_ (.A1(_3425_),
    .A2(_3721_),
    .B1(_3722_),
    .B2(_3391_),
    .ZN(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8420_ (.A1(_2544_),
    .A2(_3715_),
    .B(_3723_),
    .C(_3155_),
    .ZN(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8421_ (.A1(_3563_),
    .A2(_3718_),
    .ZN(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8422_ (.A1(_2261_),
    .A2(_2481_),
    .B(_3725_),
    .ZN(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8423_ (.A1(_1221_),
    .A2(_3647_),
    .B1(_3726_),
    .B2(_2371_),
    .C(_3106_),
    .ZN(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8424_ (.A1(_1221_),
    .A2(_3421_),
    .B(_3388_),
    .ZN(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8425_ (.A1(_2353_),
    .A2(_3724_),
    .B1(_3727_),
    .B2(_2496_),
    .C(_3728_),
    .ZN(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8426_ (.A1(net40),
    .A2(_3418_),
    .B(_2402_),
    .ZN(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8427_ (.A1(_3729_),
    .A2(_3730_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8428_ (.A1(_4034_),
    .A2(_1397_),
    .ZN(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8429_ (.I(_3731_),
    .Z(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8430_ (.I(_3732_),
    .Z(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8431_ (.I(_3731_),
    .ZN(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8432_ (.A1(_4186_),
    .A2(_4198_),
    .A3(_3734_),
    .ZN(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8433_ (.I(_3735_),
    .Z(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8434_ (.A1(\as2650.r123[2][0] ),
    .A2(_3736_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8435_ (.I(_4199_),
    .Z(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8436_ (.A1(_3738_),
    .A2(_1804_),
    .ZN(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8437_ (.A1(_4185_),
    .A2(_3733_),
    .B(_3737_),
    .C(_3739_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8438_ (.A1(_3738_),
    .A2(_1897_),
    .ZN(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8439_ (.I(_3735_),
    .Z(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8440_ (.A1(\as2650.r123[2][1] ),
    .A2(_3741_),
    .ZN(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8441_ (.A1(_0303_),
    .A2(_3733_),
    .B(_3740_),
    .C(_3742_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8442_ (.A1(_3738_),
    .A2(_1946_),
    .ZN(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8443_ (.A1(\as2650.r123[2][2] ),
    .A2(_3741_),
    .ZN(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8444_ (.A1(_0396_),
    .A2(_3733_),
    .B(_3743_),
    .C(_3744_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8445_ (.A1(_3738_),
    .A2(_1989_),
    .ZN(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8446_ (.A1(\as2650.r123[2][3] ),
    .A2(_3741_),
    .ZN(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8447_ (.A1(_0493_),
    .A2(_3733_),
    .B(_3745_),
    .C(_3746_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8448_ (.A1(_4217_),
    .A2(_2029_),
    .ZN(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8449_ (.A1(\as2650.r123[2][4] ),
    .A2(_3741_),
    .ZN(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8450_ (.A1(_0599_),
    .A2(_3732_),
    .B(_3747_),
    .C(_3748_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8451_ (.A1(_4217_),
    .A2(_2058_),
    .ZN(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8452_ (.A1(\as2650.r123[2][5] ),
    .A2(_3736_),
    .ZN(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8453_ (.A1(_0687_),
    .A2(_3732_),
    .B(_3749_),
    .C(_3750_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8454_ (.A1(\as2650.r123[2][6] ),
    .A2(_3736_),
    .ZN(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8455_ (.A1(_0496_),
    .A2(_2082_),
    .B1(_3732_),
    .B2(_0771_),
    .C(_3751_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8456_ (.A1(_0890_),
    .A2(_3734_),
    .B1(_3736_),
    .B2(\as2650.r123[2][7] ),
    .ZN(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8457_ (.A1(_0496_),
    .A2(_2103_),
    .B(_3752_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8458_ (.A1(_2258_),
    .A2(_1726_),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8459_ (.A1(_2470_),
    .A2(_1727_),
    .B(_3753_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8460_ (.I(_1535_),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8461_ (.A1(_3754_),
    .A2(_1726_),
    .ZN(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8462_ (.A1(_2459_),
    .A2(_1727_),
    .B(_3755_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8463_ (.I(_3174_),
    .Z(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8464_ (.A1(_2992_),
    .A2(_1384_),
    .ZN(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _8465_ (.A1(_0438_),
    .A2(_1410_),
    .A3(_2497_),
    .A4(_2369_),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8466_ (.A1(_2170_),
    .A2(_2584_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8467_ (.A1(_1596_),
    .A2(_3759_),
    .ZN(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8468_ (.A1(_1064_),
    .A2(_3164_),
    .B(_1555_),
    .ZN(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8469_ (.A1(_1412_),
    .A2(_1273_),
    .B(_1733_),
    .C(_1280_),
    .ZN(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8470_ (.A1(_1419_),
    .A2(_3762_),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8471_ (.A1(_4164_),
    .A2(_4194_),
    .B1(_1102_),
    .B2(_1101_),
    .C(_1254_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8472_ (.A1(_2466_),
    .A2(_3764_),
    .B(_2328_),
    .C(_3131_),
    .ZN(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8473_ (.A1(_1392_),
    .A2(_2368_),
    .A3(_3763_),
    .A4(_3765_),
    .ZN(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8474_ (.A1(_3758_),
    .A2(_3760_),
    .A3(_3761_),
    .A4(_3766_),
    .ZN(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8475_ (.A1(_1411_),
    .A2(_1579_),
    .ZN(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8476_ (.I(_1402_),
    .ZN(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8477_ (.A1(_2361_),
    .A2(_1092_),
    .B1(_1262_),
    .B2(_3769_),
    .C(_2594_),
    .ZN(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8478_ (.A1(_2601_),
    .A2(_3768_),
    .A3(_3770_),
    .ZN(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8479_ (.A1(_3757_),
    .A2(_3767_),
    .A3(_3771_),
    .ZN(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8480_ (.A1(_1725_),
    .A2(_3756_),
    .B(_3772_),
    .ZN(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8481_ (.A1(_2354_),
    .A2(_1432_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8482_ (.A1(_0992_),
    .A2(_2398_),
    .B1(_3774_),
    .B2(_1725_),
    .ZN(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8483_ (.A1(_1063_),
    .A2(_0967_),
    .Z(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8484_ (.A1(_0973_),
    .A2(_2977_),
    .B1(_3776_),
    .B2(_2302_),
    .ZN(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8485_ (.A1(_3070_),
    .A2(_3775_),
    .B(_3777_),
    .ZN(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8486_ (.A1(_3773_),
    .A2(_3778_),
    .ZN(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8487_ (.A1(_1063_),
    .A2(_3773_),
    .B(_3779_),
    .C(_3624_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8488_ (.A1(_1531_),
    .A2(_3756_),
    .B(_3772_),
    .ZN(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8489_ (.A1(_2576_),
    .A2(_2429_),
    .B(_2430_),
    .C(_1425_),
    .ZN(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8490_ (.A1(_2695_),
    .A2(_1593_),
    .ZN(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8491_ (.A1(_3781_),
    .A2(_3782_),
    .B(_2528_),
    .ZN(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8492_ (.A1(_2528_),
    .A2(_0927_),
    .B(_3783_),
    .ZN(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8493_ (.A1(_0978_),
    .A2(_3780_),
    .B1(_3784_),
    .B2(_3772_),
    .ZN(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8494_ (.A1(_3242_),
    .A2(_3785_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8495_ (.A1(_1717_),
    .A2(_3756_),
    .B(_3772_),
    .ZN(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8496_ (.A1(_2576_),
    .A2(_2425_),
    .B(_3070_),
    .ZN(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8497_ (.A1(_0968_),
    .A2(_3070_),
    .B1(_2426_),
    .B2(_3787_),
    .C(_3786_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8498_ (.A1(_0968_),
    .A2(_3786_),
    .B(_3788_),
    .C(_3624_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8499_ (.I(_0439_),
    .Z(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8500_ (.I(_1418_),
    .Z(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8501_ (.A1(_3790_),
    .A2(_1426_),
    .B(_3789_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8502_ (.A1(_3789_),
    .A2(_0544_),
    .B1(_2446_),
    .B2(_3791_),
    .ZN(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8503_ (.A1(_3266_),
    .A2(_3792_),
    .B(_3288_),
    .ZN(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8504_ (.A1(_2280_),
    .A2(_3793_),
    .ZN(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8505_ (.A1(_1570_),
    .A2(_1431_),
    .A3(_2473_),
    .ZN(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8506_ (.A1(_1428_),
    .A2(_3795_),
    .ZN(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8507_ (.A1(_1320_),
    .A2(_1582_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8508_ (.A1(_1247_),
    .A2(_2591_),
    .A3(_1420_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8509_ (.A1(_0473_),
    .A2(_4279_),
    .B(_3798_),
    .ZN(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8510_ (.A1(_1591_),
    .A2(_1417_),
    .A3(_3175_),
    .ZN(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _8511_ (.A1(_1265_),
    .A2(_3797_),
    .A3(_3799_),
    .A4(_3800_),
    .Z(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8512_ (.A1(_3760_),
    .A2(_3801_),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8513_ (.A1(_1590_),
    .A2(_3802_),
    .ZN(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8514_ (.A1(_1841_),
    .A2(_2992_),
    .B1(_2375_),
    .B2(_3756_),
    .ZN(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8515_ (.A1(_3789_),
    .A2(_3804_),
    .ZN(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8516_ (.A1(_1720_),
    .A2(_2299_),
    .ZN(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8517_ (.A1(_1841_),
    .A2(_2273_),
    .B(_1566_),
    .C(_2301_),
    .ZN(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8518_ (.A1(_1392_),
    .A2(_2381_),
    .A3(_3806_),
    .A4(_3807_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8519_ (.A1(_3761_),
    .A2(_3803_),
    .A3(_3805_),
    .A4(_3808_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8520_ (.A1(_2459_),
    .A2(_0548_),
    .B(_3796_),
    .C(_3809_),
    .ZN(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8521_ (.A1(_3796_),
    .A2(_3809_),
    .ZN(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8522_ (.A1(\as2650.psl[5] ),
    .A2(_3811_),
    .ZN(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8523_ (.A1(_3794_),
    .A2(_3810_),
    .B(_3812_),
    .C(_3624_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8524_ (.A1(_0747_),
    .A2(_1518_),
    .ZN(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8525_ (.A1(_0850_),
    .A2(_1345_),
    .ZN(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8526_ (.A1(_0462_),
    .A2(_0850_),
    .B(_3814_),
    .ZN(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8527_ (.A1(_3815_),
    .A2(_0492_),
    .ZN(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8528_ (.A1(_4169_),
    .A2(_4182_),
    .B(_0300_),
    .ZN(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8529_ (.A1(_4169_),
    .A2(_4182_),
    .A3(_0299_),
    .ZN(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8530_ (.A1(_0348_),
    .A2(_0478_),
    .B1(_3817_),
    .B2(_4289_),
    .C(_3818_),
    .ZN(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8531_ (.A1(_0349_),
    .A2(_0478_),
    .ZN(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8532_ (.A1(_3816_),
    .A2(_3819_),
    .A3(_3820_),
    .ZN(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8533_ (.A1(_3815_),
    .A2(_0491_),
    .B1(_0539_),
    .B2(_0547_),
    .ZN(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8534_ (.I(_3822_),
    .ZN(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8535_ (.A1(_0539_),
    .A2(_0547_),
    .B1(_3821_),
    .B2(_3823_),
    .ZN(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8536_ (.A1(_0648_),
    .A2(_0759_),
    .ZN(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8537_ (.A1(_0648_),
    .A2(_0759_),
    .ZN(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8538_ (.A1(_0747_),
    .A2(_1518_),
    .B1(_3824_),
    .B2(_3825_),
    .C(_3826_),
    .ZN(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8539_ (.A1(_0862_),
    .A2(_1514_),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8540_ (.A1(_3813_),
    .A2(_3827_),
    .B(_3828_),
    .ZN(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8541_ (.A1(_0862_),
    .A2(_1514_),
    .ZN(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8542_ (.A1(_1571_),
    .A2(_3830_),
    .ZN(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8543_ (.A1(_2323_),
    .A2(_3790_),
    .ZN(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8544_ (.A1(_4214_),
    .A2(_2354_),
    .B1(_3832_),
    .B2(_1530_),
    .C(_1561_),
    .ZN(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8545_ (.A1(_3789_),
    .A2(_1624_),
    .B(_3833_),
    .ZN(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8546_ (.A1(_3266_),
    .A2(_4251_),
    .ZN(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8547_ (.A1(_3266_),
    .A2(_3834_),
    .B(_3835_),
    .C(_2279_),
    .ZN(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8548_ (.A1(_1717_),
    .A2(_3795_),
    .ZN(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8549_ (.A1(_3809_),
    .A2(_3837_),
    .ZN(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8550_ (.A1(_3836_),
    .A2(_3838_),
    .ZN(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8551_ (.A1(_3829_),
    .A2(_3831_),
    .B(_3839_),
    .ZN(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8552_ (.A1(\as2650.carry ),
    .A2(_3838_),
    .B(_2402_),
    .ZN(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8553_ (.A1(_3840_),
    .A2(_3841_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8554_ (.A1(_1379_),
    .A2(_1382_),
    .ZN(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8555_ (.A1(_2279_),
    .A2(_2255_),
    .A3(_1431_),
    .ZN(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _8556_ (.A1(_1414_),
    .A2(_2523_),
    .B(_2287_),
    .C(_2231_),
    .ZN(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8557_ (.A1(_3842_),
    .A2(_3803_),
    .A3(_3843_),
    .A4(_3844_),
    .ZN(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8558_ (.A1(_3790_),
    .A2(_2434_),
    .B(_2432_),
    .ZN(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8559_ (.A1(_2280_),
    .A2(_3846_),
    .B(_3845_),
    .ZN(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8560_ (.A1(_0861_),
    .A2(_1514_),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8561_ (.A1(_3848_),
    .A2(_3830_),
    .B(_1688_),
    .C(_1502_),
    .ZN(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8562_ (.A1(_3230_),
    .A2(_3845_),
    .B1(_3847_),
    .B2(_3849_),
    .C(_2493_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8563_ (.A1(_3754_),
    .A2(_2442_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8564_ (.A1(_2635_),
    .A2(_1406_),
    .B(_2319_),
    .ZN(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8565_ (.A1(_4202_),
    .A2(_2323_),
    .ZN(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8566_ (.A1(_1378_),
    .A2(_1396_),
    .A3(_3851_),
    .A4(_3852_),
    .ZN(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8567_ (.A1(_1393_),
    .A2(_1589_),
    .A3(_3853_),
    .ZN(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8568_ (.I(_3854_),
    .Z(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8569_ (.A1(_3850_),
    .A2(_3855_),
    .B(_4036_),
    .ZN(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8570_ (.A1(_1350_),
    .A2(_2437_),
    .B1(_3832_),
    .B2(_3754_),
    .ZN(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8571_ (.A1(_3855_),
    .A2(_3857_),
    .Z(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8572_ (.A1(_3856_),
    .A2(_3858_),
    .B(_2492_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8573_ (.A1(_3246_),
    .A2(_2442_),
    .ZN(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8574_ (.A1(_3855_),
    .A2(_3859_),
    .B(_1841_),
    .ZN(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8575_ (.A1(_1344_),
    .A2(_2437_),
    .B1(_3832_),
    .B2(_3246_),
    .ZN(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8576_ (.A1(_3855_),
    .A2(_3861_),
    .Z(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8577_ (.A1(_3860_),
    .A2(_3862_),
    .B(_2492_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8578_ (.A1(_2251_),
    .A2(_2433_),
    .B(_3854_),
    .ZN(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8579_ (.A1(\as2650.psl[1] ),
    .A2(_3863_),
    .ZN(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8580_ (.A1(_3790_),
    .A2(_2429_),
    .B(_2430_),
    .C(_3863_),
    .ZN(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8581_ (.A1(_1635_),
    .A2(_3865_),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8582_ (.A1(_3864_),
    .A2(_3866_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8583_ (.I(net27),
    .ZN(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8584_ (.A1(_3885_),
    .A2(_2329_),
    .A3(_3761_),
    .ZN(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _8585_ (.A1(_4191_),
    .A2(_1383_),
    .A3(_3851_),
    .A4(_3868_),
    .ZN(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8586_ (.I(_3869_),
    .Z(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8587_ (.A1(_1739_),
    .A2(_2441_),
    .B(_3870_),
    .ZN(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8588_ (.A1(_1739_),
    .A2(_2433_),
    .A3(_2576_),
    .ZN(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8589_ (.A1(_1167_),
    .A2(_2436_),
    .B(_3872_),
    .ZN(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8590_ (.A1(_3867_),
    .A2(_3871_),
    .B1(_3873_),
    .B2(_3870_),
    .C(_2493_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8591_ (.A1(_3754_),
    .A2(_2441_),
    .B(_3869_),
    .ZN(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8592_ (.A1(_1025_),
    .A2(_2355_),
    .B1(_3774_),
    .B2(_1535_),
    .ZN(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8593_ (.I(_3875_),
    .ZN(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8594_ (.A1(\as2650.psu[4] ),
    .A2(_3874_),
    .B1(_3876_),
    .B2(_3870_),
    .ZN(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8595_ (.A1(_3242_),
    .A2(_3877_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8596_ (.A1(_2258_),
    .A2(_2441_),
    .B(_3869_),
    .ZN(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8597_ (.A1(_1005_),
    .A2(_2355_),
    .B1(_3774_),
    .B2(_3246_),
    .ZN(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8598_ (.I(_3879_),
    .ZN(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8599_ (.A1(\as2650.psu[3] ),
    .A2(_3878_),
    .B1(_3880_),
    .B2(_3870_),
    .ZN(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8600_ (.A1(_2492_),
    .A2(_3881_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8601_ (.D(_0000_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8602_ (.D(_0001_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8603_ (.D(_0002_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8604_ (.D(_0003_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8605_ (.D(_0004_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8606_ (.D(_0005_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8607_ (.D(_0006_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8608_ (.D(_0007_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8609_ (.D(_0008_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8610_ (.D(_0009_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8611_ (.D(_0010_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8612_ (.D(_0011_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8613_ (.D(_0012_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8614_ (.D(_0013_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8615_ (.D(_0014_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8616_ (.D(_0015_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8617_ (.D(_0016_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8618_ (.D(_0017_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8619_ (.D(_0018_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8620_ (.D(_0019_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8621_ (.D(_0020_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8622_ (.D(_0021_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8623_ (.D(_0022_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8624_ (.D(_0023_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8625_ (.D(_0024_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8626_ (.D(_0025_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8627_ (.D(_0026_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8628_ (.D(_0027_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8629_ (.D(_0028_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8630_ (.D(_0029_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8631_ (.D(_0030_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8632_ (.D(_0031_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8633_ (.D(_0032_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8634_ (.D(_0033_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8635_ (.D(_0034_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8636_ (.D(_0035_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8637_ (.D(_0036_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8638_ (.D(_0037_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8639_ (.D(_0038_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8640_ (.D(_0039_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8641_ (.D(_0040_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\as2650.r123_2[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8642_ (.D(_0041_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\as2650.r123_2[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8643_ (.D(_0042_),
    .CLK(clknet_opt_2_1_wb_clk_i),
    .Q(\as2650.r123_2[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8644_ (.D(_0043_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.r123_2[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8645_ (.D(_0044_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.r123_2[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8646_ (.D(_0045_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8647_ (.D(_0046_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123_2[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8648_ (.D(_0047_),
    .CLK(clknet_opt_3_0_wb_clk_i),
    .Q(\as2650.r123_2[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8649_ (.D(_0048_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8650_ (.D(_0049_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8651_ (.D(_0050_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8652_ (.D(_0051_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8653_ (.D(_0052_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8654_ (.D(_0053_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8655_ (.D(_0054_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8656_ (.D(_0055_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8657_ (.D(_0056_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8658_ (.D(_0057_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8659_ (.D(_0058_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8660_ (.D(_0059_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8661_ (.D(_0060_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8662_ (.D(_0061_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8663_ (.D(_0062_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8664_ (.D(_0063_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8665_ (.D(_0064_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8666_ (.D(_0065_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8667_ (.D(_0066_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8668_ (.D(_0067_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8669_ (.D(_0068_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8670_ (.D(_0069_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8671_ (.D(_0070_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8672_ (.D(_0071_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8673_ (.D(_0072_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8674_ (.D(_0073_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8675_ (.D(_0074_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8676_ (.D(_0075_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8677_ (.D(_0076_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8678_ (.D(_0077_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8679_ (.D(_0078_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8680_ (.D(_0079_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8681_ (.D(_0080_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8682_ (.D(_0081_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8683_ (.D(_0082_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8684_ (.D(_0083_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8685_ (.D(_0084_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8686_ (.D(_0085_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8687_ (.D(_0086_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8688_ (.D(_0087_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8689_ (.D(_0088_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8690_ (.D(_0089_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8691_ (.D(_0090_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8692_ (.D(_0091_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8693_ (.D(_0092_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8694_ (.D(_0093_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8695_ (.D(_0094_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8696_ (.D(_0095_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8697_ (.D(_0096_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8698_ (.D(_0097_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8699_ (.D(_0098_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8700_ (.D(_0099_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8701_ (.D(_0100_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8702_ (.D(_0101_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8703_ (.D(_0102_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8704_ (.D(_0103_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8705_ (.D(_0104_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8706_ (.D(_0105_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8707_ (.D(_0106_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8708_ (.D(_0107_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8709_ (.D(_0108_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8710_ (.D(_0109_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8711_ (.D(_0110_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8712_ (.D(_0111_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8713_ (.D(_0112_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8714_ (.D(_0113_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8715_ (.D(_0114_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8716_ (.D(_0115_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8717_ (.D(_0116_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8718_ (.D(_0117_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8719_ (.D(_0118_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8720_ (.D(_0119_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8721_ (.D(_0120_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8722_ (.D(_0121_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8723_ (.D(_0122_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8724_ (.D(_0123_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8725_ (.D(_0124_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8726_ (.D(_0125_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8727_ (.D(_0126_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8728_ (.D(_0127_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8729_ (.D(_0128_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8730_ (.D(_0129_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8731_ (.D(_0130_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8732_ (.D(_0131_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8733_ (.D(_0132_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8734_ (.D(_0133_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8735_ (.D(_0134_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8736_ (.D(_0135_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8737_ (.D(_0136_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8738_ (.D(_0137_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8739_ (.D(_0138_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8740_ (.D(_0139_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8741_ (.D(_0140_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8742_ (.D(_0141_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8743_ (.D(_0142_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8744_ (.D(_0143_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8745_ (.D(_0144_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8746_ (.D(_0145_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8747_ (.D(_0146_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8748_ (.D(_0147_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8749_ (.D(_0148_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8750_ (.D(_0149_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8751_ (.D(_0150_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8752_ (.D(_0151_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8753_ (.D(_0152_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8754_ (.D(_0153_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8755_ (.D(_0154_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8756_ (.D(_0155_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8757_ (.D(_0156_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8758_ (.D(_0157_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8759_ (.D(_0158_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8760_ (.D(_0159_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8761_ (.D(_0160_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8762_ (.D(_0161_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8763_ (.D(_0162_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8764_ (.D(_0163_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8765_ (.D(_0164_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8766_ (.D(_0165_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8767_ (.D(_0166_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8768_ (.D(_0167_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8769_ (.D(_0168_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _8770_ (.D(_0169_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8771_ (.D(_0170_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8772_ (.D(_0171_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8773_ (.D(_0172_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8774_ (.D(_0173_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8775_ (.D(_0174_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8776_ (.D(_0175_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8777_ (.D(_0176_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8778_ (.D(_0177_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8779_ (.D(_0178_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8780_ (.D(_0179_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8781_ (.D(_0180_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8782_ (.D(_0181_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8783_ (.D(_0182_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8784_ (.D(_0183_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8785_ (.D(_0184_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8786_ (.D(_0185_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _8787_ (.D(_0186_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _8788_ (.D(_0187_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8789_ (.D(_0188_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8790_ (.D(_0189_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8791_ (.D(_0190_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8792_ (.D(_0191_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8793_ (.D(_0192_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8794_ (.D(_0193_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8795_ (.D(_0194_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8796_ (.D(_0195_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8797_ (.D(_0196_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8798_ (.D(_0197_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8799_ (.D(_0198_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8800_ (.D(_0199_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8801_ (.D(_0200_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8802_ (.D(_0201_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8803_ (.D(_0202_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8804_ (.D(_0203_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8805_ (.D(_0204_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8806_ (.D(_0205_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8807_ (.D(_0206_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8808_ (.D(_0207_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8809_ (.D(_0208_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8810_ (.D(_0209_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8811_ (.D(_0210_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8812_ (.D(_0211_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8813_ (.D(_0212_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8814_ (.D(_0213_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8815_ (.D(_0214_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8816_ (.D(_0215_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8817_ (.D(_0216_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8818_ (.D(_0217_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8819_ (.D(_0218_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8820_ (.D(_0219_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8821_ (.D(_0220_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8822_ (.D(_0221_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8823_ (.D(_0222_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8824_ (.D(_0223_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8825_ (.D(_0224_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8826_ (.D(_0225_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8827_ (.D(_0226_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8828_ (.D(_0227_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8829_ (.D(_0228_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8830_ (.D(_0229_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8831_ (.D(_0230_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8832_ (.D(_0231_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8833_ (.D(_0232_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8834_ (.D(_0233_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8835_ (.D(_0234_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8836_ (.D(_0235_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8837_ (.D(_0236_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8838_ (.D(_0237_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8839_ (.D(_0238_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8840_ (.D(_0239_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8841_ (.D(_0240_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8842_ (.D(_0241_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8843_ (.D(_0242_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8844_ (.D(_0243_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8845_ (.D(_0244_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8846_ (.D(_0245_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8847_ (.D(_0246_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8848_ (.D(_0247_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8849_ (.D(_0248_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8850_ (.D(_0249_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8851_ (.D(_0250_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8852_ (.D(_0251_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8853_ (.D(_0252_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8854_ (.D(_0253_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8855_ (.D(_0254_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8856_ (.D(_0255_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8857_ (.D(_0256_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8858_ (.D(_0257_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8859_ (.D(_0258_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8860_ (.D(_0259_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8861_ (.D(_0260_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8862_ (.D(_0261_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8863_ (.D(_0262_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8864_ (.D(_0263_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8865_ (.D(_0264_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8866_ (.D(_0265_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8867_ (.D(_0266_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8868_ (.D(_0267_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8869_ (.D(_0268_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8870_ (.D(_0269_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8871_ (.D(_0270_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8872_ (.D(_0271_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8873_ (.D(_0272_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8874_ (.D(_0273_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8875_ (.D(_0274_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8876_ (.D(_0275_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8877_ (.D(_0276_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8878_ (.D(_0277_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8879_ (.D(_0278_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8880_ (.D(_0279_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8881_ (.D(_0280_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8882_ (.D(_0281_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8883_ (.D(_0282_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8884_ (.D(_0283_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_89 (.Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_90 (.Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_91 (.Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_92 (.Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_93 (.Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_88 (.Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8926_ (.I(net46),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8927_ (.I(net46),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8928_ (.I(net47),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8929_ (.I(net46),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8930_ (.I(net47),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8931_ (.I(net47),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8932_ (.I(net46),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(io_in[5]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input6 (.I(io_in[6]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input7 (.I(io_in[7]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(io_in[8]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(io_in[9]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(wb_rst_i),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net49),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net52),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net13),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout50 (.I(net37),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout51 (.I(net33),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net29),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_opt_1_1_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_1_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_opt_1_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_1_wb_clk_i (.I(clknet_opt_2_0_wb_clk_i),
    .Z(clknet_opt_2_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_3_0_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__D (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8762__D (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__D (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__D (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__D (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8791__D (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__D (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__D (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__D (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__D (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__D (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8879__D (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__C (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__I (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A3 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A3 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A3 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__I (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__B1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A4 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__B2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__I (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__B (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__I (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__B (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__B2 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A2 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__B2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__B2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__B2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__B2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__B2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__I (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__B2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__B1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__B1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A4 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__I (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A4 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A3 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A3 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__I (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__I (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__B (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__B2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A3 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__I (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__B (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__B (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A3 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__I (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A4 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A4 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__B1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__I (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__I (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__S (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__S (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__S (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__B2 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__I (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__I (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A3 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__B2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__I (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__I (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__I (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__B1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__I (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__I (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__I (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__I (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__B (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__I (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__I (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__B (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A4 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__C (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__C (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__B1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__B1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A3 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A3 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__S (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__B (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__B (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__I (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__B (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__C (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__B (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__B (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__B1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__B2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__B2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A4 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A4 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__I (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A3 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A2 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__I (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__B2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__B1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__B2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__B (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8535__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__B1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A4 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8535__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__B2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A3 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__I (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__I (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__I (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__I (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__I (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__I (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A3 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__B1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A3 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__I (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__I (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__A1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__B1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A3 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__B2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__B2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__I (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__I (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__I (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__I (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__B (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A4 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__I (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__B1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__B1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__B1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__B (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__B (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A3 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__I (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__C1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__B1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__I (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__I (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__I (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__B1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__C2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__I (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__I (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__B2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__B2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__B1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__I (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__I (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__I (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A3 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A3 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A3 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__I (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__B1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A3 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__B (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__B1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A1 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__A2 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__B2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__B1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__I (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__B1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__I (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__I (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__I (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__I (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__B (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__C (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__B2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A3 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__I0 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__I (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__B2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A4 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__I (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__I (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A3 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__B1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__I (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A3 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A3 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__I (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A2 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__B1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A4 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A3 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__B (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__I (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__I (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__I (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__B2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__B1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__B (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__B1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A4 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A4 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A3 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__C (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A1 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A1 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__I (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A3 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A3 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A3 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A3 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A3 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A3 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A2 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__B1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__I (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__S0 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__C1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__S1 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__I (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__A1 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__B2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__B2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__I (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__I (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__B2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__B2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__B1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__I (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__B1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__B1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__B1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__S (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__S (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__I (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__S0 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__S (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__S0 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__S (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__B2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__I (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__B (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__B (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__B (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__B (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__B2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__B2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__I (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__B2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__B2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__B2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__B2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__B2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__B2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__B2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__I (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__I (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__I (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__I (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__B2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__B2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__B2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__B2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__I (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__I (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__C (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__C (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__I (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__C (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__C (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__C (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__C (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__B2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__A1 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__B1 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__I (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__B2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__I (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__I (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__I (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__A2 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__B2 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__B2 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__B2 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__C (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__C (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__C (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__I (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__B2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__C (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__C (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__I (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__C (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__C (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__C (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__C (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__C (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__C (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__I (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__A1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__S1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__S1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__B1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A3 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__I (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__B1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__B1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__C (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__B2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__B2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__I (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__B2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__B2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__B2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__S0 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__S0 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__S0 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__S1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__S1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__S1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__A2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__B1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__B2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__B1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__C (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__I (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__B2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__B1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__B1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__C (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__I (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__B1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__B1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__C (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__B2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__B (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__B (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__B (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__I (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A2 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__I (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__I (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__I (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A3 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__S (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__S (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__B (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__I (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__I (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A3 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__I (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__B (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__I (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__I (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__I (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__I (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__I (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__B (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__I (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__I (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A3 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__B (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__B (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__B2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__B2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__B1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__B (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__I (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__I (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A3 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__B (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__I (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__I (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A1 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__C (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__C (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A3 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__A2 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__A2 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__I (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__I (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__I (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__I (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__I1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__I (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__I (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A2 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A2 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__I (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__I (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A3 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__I (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__I (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__I (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__B (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__I (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__I (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__B2 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__I (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__I (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A1 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__I (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__I (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__I (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A2 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__I (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__B (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__I (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__I0 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__I0 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A1 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__A1 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__A1 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__I1 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__I (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__I (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__I (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__I (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__I (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__I (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__I (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__I (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__I (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__I (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__I (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__I (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__I (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__B2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__I (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A3 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A3 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__I (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A4 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__I (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__I (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__B (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__B (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A3 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__I (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__I (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__I (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__C (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__I (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__I (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__I (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__B (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A3 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__I (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__B1 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__I (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A1 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A3 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A3 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__C (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7751__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__I (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__I (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__I (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__I (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__I (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__I (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__B (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__I (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__B1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__I (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__B2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__C (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__I (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__I (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__I (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A3 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A3 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__I (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A1 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A4 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A4 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__I (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__I (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A3 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A3 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__I (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__B (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__I (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__I (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__B1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__I (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A1 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__I (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__C (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__I (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__B (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__B2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__I (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__I (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__B2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__B (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__I (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__C (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A3 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A2 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A3 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__B (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__I (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__I (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A4 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__A2 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A2 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A3 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__I (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__I (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__I (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__I (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__B2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__B2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A2 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A2 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__I (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__B (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__I (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__B (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__I (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__I (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A2 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A4 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__I (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A3 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__I (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A1 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A3 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A2 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A3 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A4 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A3 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__I (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__I (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__I (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__B (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__C (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__B (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A3 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__C (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__A1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A2 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A3 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A3 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A2 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__I (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A3 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A3 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__I (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A3 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__I (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__I (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__A1 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__I (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__C (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A3 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__I (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__C (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__C (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__B (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A3 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A3 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__C (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__A1 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A2 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A4 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A3 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__B (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__C (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__B (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__A1 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__I (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A2 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__B (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__I (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__B (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__I (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__B2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__B (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__I (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A3 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__B (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__C (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__C (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__C (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__C (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__I (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__I (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A2 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A2 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A2 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A2 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__I (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__I (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__I (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__I (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A2 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A2 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A2 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A2 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A2 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__I (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__I (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__I (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__I (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__I (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A2 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A2 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A2 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__I (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__I (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__I (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__I (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__I (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__I (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__C (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__B (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__B (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A3 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__A2 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__A2 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__A2 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__C (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__C (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__B (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__B (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__I (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__I (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__C (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__I (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__I (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__B2 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A3 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__I (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__I (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A4 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__B2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7677__A2 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__B (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__A2 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__I (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__C1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__I (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__I (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__I (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__I (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A3 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A1 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__A1 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__B (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__I (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__C (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__C (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__C (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__B (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__B (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__I (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__C (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__B (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__C (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__B (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__C (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__B (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__B (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A1 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__C (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__B (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__B (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__I (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__B2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__C (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__C (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__B (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__B1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__B (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__B1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__B (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A2 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A4 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__A2 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__A2 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__B (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__I (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__I (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A3 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A2 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A3 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__B1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__I (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__B2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A3 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A3 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A2 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A3 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__B (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__C (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A3 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__B (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A4 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A2 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__I (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__A3 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__I (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A2 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A3 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A3 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A3 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__C (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A4 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__S (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A3 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__B1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__B2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__I (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__B1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A2 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__B1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__B2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A3 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A2 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A3 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__B (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__B (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__A2 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__B (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__C (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__I0 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__C (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__I (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__I (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A2 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A1 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A1 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A1 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A2 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A3 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__B (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__B1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__I (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__B1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__I (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A2 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A2 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__B (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__B1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__C (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__A1 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__B2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__C2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__C (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__B2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__C (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__B2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__B (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__C (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__I (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__C (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__I (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__I (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__B (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__C (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__B (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__C (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__C (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__I1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A2 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A3 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__B1 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__B1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__B1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__B (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__B (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__A1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__I (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A1 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__B2 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__A2 (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A2 (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A2 (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A2 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__B2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__B2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A3 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__I (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__I (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__B (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__I (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__I (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__I (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__I (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__C (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7562__C (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__I (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__I (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__B2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A2 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A2 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A2 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A2 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__I (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__I (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__I (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__I (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__I (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__I (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A3 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__I (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__A1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__I (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A3 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A2 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A3 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A1 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A1 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A3 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__C (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__I (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__I (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__C (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__C (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__I (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A3 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A4 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A3 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__B (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A3 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__I (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__I (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__B (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__B (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A3 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A2 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A2 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A2 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A2 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__S (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__I (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__B (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A4 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__I (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A4 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A3 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A3 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A2 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A2 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A2 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__I (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__I (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__I (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__I (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A3 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__C (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__A2 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A2 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A2 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A2 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__C (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__I (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__B (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__I (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__I (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__B (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__I (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__B (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__I (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__B (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A2 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__B1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__B1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__B2 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__C (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__B (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__C (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__C (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__C (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A2 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__B1 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A2 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__A2 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A2 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__B1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__A1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__B1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A1 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__I (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__A2 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A2 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A1 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A1 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__B (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A1 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A1 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__I (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A1 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A1 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__B (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__C (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__C (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A1 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A2 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__A1 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__B1 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__I (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__B1 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__A1 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__C (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A2 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A2 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__B1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A2 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A1 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A3 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A2 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A2 (.I(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A2 (.I(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__A1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__A1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A2 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A2 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A2 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A2 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A2 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A2 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__I (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__B (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__C (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__A2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A3 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__I (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__C (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__A2 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A2 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__A2 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A2 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__A2 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__A2 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__B1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__A2 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__A2 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__I (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__I (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__A2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A2 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A2 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A2 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A2 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__C (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__I (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__I (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__I (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__A1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__B1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__I (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A1 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__I (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__C (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__A3 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__B1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__B1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__B1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__B1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__B (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A3 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__B1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__B1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__B1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__B1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A1 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__B (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__I (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A2 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A1 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__A2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__C (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__C (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__I (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__I (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A3 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A3 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A2 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A2 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A4 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A3 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__B (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__C (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__A2 (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A2 (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__I (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A1 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A2 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__I (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A1 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__C (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__I (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__I (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__B1 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__C (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__I (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A2 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__B2 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A2 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__A3 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__B1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A3 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A4 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A2 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A3 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A2 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A1 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A3 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A3 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A3 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A4 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__A1 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A3 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__A4 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A3 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__A2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__S (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__I (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__A1 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A1 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__A1 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A1 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A1 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__A1 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A1 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A1 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A2 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A2 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A2 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__A2 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A2 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__I0 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__I (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__I1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__B (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A2 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__I1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__B2 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__C2 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__I (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A1 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__I (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__B2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A4 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__B (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__A1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A1 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__C (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__B2 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__I (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__B2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__C (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__I (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__I (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__I (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__A1 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A2 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__B (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__B (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__I (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A2 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A3 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__A2 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A4 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__A3 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A3 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A2 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__I (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__B2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A4 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__B1 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__A1 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A2 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__I (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A1 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__B1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A2 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__A2 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A2 (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A2 (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A2 (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A1 (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__B2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__I (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__I (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__B (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__I (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__C1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__C (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__B (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__I (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__I (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__B2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__C (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__C (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__C2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__A1 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__A1 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A1 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__B (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A2 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A4 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__B (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__B (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__I (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__B (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A3 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__A2 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A2 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__A2 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A4 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__B (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A1 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__I (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A4 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__I (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__B (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A4 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__A3 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__A1 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__I (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A3 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8070__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__A1 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A1 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__A3 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__B1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A3 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A2 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__C (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__I (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__B2 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__I (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A3 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A4 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A2 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__B (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__A2 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__A2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A2 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A2 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A2 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A3 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__A2 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__I (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__B2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__C (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A3 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__B (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__B2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__B (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__A1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A4 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A2 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A2 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A2 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__B2 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__A2 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__I (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A2 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__B1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A4 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__B1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__I (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__C (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A2 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__I (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A2 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__B (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A3 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__B2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__B2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__B (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A4 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A2 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A2 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A2 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A3 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A2 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__I (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__C (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__B (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__B2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A3 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__I (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__I (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__C (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__C (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__B (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__B (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A2 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A3 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__A2 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__I (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A2 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A2 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A2 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__C (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__B (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A2 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A2 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__B (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__B (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8426__B (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__B (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__B (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A3 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__B (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__I (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__I (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__I (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__I (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A2 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__A3 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__B (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__B (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__I (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__I (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__I (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__I (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__C (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__C (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__C (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__C (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__I (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__I (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__S (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__S (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__S (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__I (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A2 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A2 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A2 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A1 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A2 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A2 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A1 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__C (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__I (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__I (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__B (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__B1 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A2 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__B2 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__I (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A2 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__A2 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__A2 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A3 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__B (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__B (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A4 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__B (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__B (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A3 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__B (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__A2 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__S (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A2 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A2 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A1 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A2 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__A2 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__A2 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__A2 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A2 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__A2 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__A2 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A1 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A2 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__I0 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__B1 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__I0 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__B (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__A1 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A1 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__A1 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A1 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__C (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__C (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__C (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__I (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__C (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A1 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A1 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A1 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A4 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A1 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__I (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A1 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A1 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A1 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A2 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__A2 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A2 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__I (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A2 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A1 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__I (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__I (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A2 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__B2 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__B (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__B (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A1 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A1 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__I (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__C (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__B (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__B2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__C (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A1 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__A1 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__C (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A1 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__I (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__I (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A3 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A3 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__B2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__B (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__B (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A1 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__B (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__B1 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__I (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__B (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A3 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__I (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__I (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A3 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__B (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__B (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__B (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__B (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__C (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__C (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__B (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__B (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__I (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__I (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__C (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__I (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__I (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__I (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__B2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A1 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A1 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A1 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A3 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__B (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__I (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__A1 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A1 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__A1 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A2 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A3 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__I (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__I (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7693__B (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A1 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__I (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__I (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__C (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A1 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A1 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A3 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__B (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__C (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__C (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__C (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A1 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__C (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A2 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__C (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__B (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A2 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A2 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A2 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__B (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__C1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__B1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__A2 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A3 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A2 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__C (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__C (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__C (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__I (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A1 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__B (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__B (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A1 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__B (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7562__A1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__A1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__C (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__B2 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__C (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__B1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__A1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A3 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A3 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__B (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__C (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__C (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__A1 (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__C (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A1 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A1 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__A1 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A2 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__B2 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A1 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__I (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__I (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A1 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A1 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A1 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A2 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__B2 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A1 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A3 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A1 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__A1 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A2 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__A1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8070__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A3 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A2 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A1 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A4 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__C (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A2 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A4 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A3 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__A1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__B1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A4 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__I (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__I (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__I (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__C (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__I (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__I (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__I (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__I (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__C (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__I (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__I (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A2 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A2 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A2 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A1 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__B2 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__A1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__A2 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__B2 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__B1 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A1 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__I (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__I (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A1 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__A1 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__B2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__B (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7641__I (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A1 (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__I (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__A1 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A1 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__I (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__I (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A2 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__B (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__A1 (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__B (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__B (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__B (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__C2 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A2 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__A1 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__C (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__B (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__I (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__A2 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__I (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__B (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__A2 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__B (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__A1 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A1 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__C2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A1 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__B1 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A2 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A2 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__I (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__I (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__I (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A2 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A2 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__B2 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__B2 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__B (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__B (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__B2 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A1 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__A1 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__I (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__I (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7602__A1 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A1 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A1 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A1 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7806__B2 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__C1 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A1 (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__I (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__I (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__I (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__C2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__A1 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__C2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__A1 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__B2 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__B2 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__B2 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__B (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__C (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__I (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__I (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__B2 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A1 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A1 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__A1 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A2 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A2 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__I (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__B (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__B (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__B (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__A1 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__B2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A1 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A1 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A1 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A2 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__B2 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__B2 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__A1 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__B2 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A1 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A1 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A1 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__A1 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A1 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A2 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__B1 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__B1 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A4 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__I (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__B1 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__I (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A1 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__A1 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__B2 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__I (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__B2 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__B (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__A1 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A3 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A2 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A1 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A1 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A1 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A3 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A4 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__B1 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__A1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__A1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__A2 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__B2 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A2 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__A2 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__A1 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A2 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A2 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A2 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A2 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__B1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__B1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__I (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__I (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__A1 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A2 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__B1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A1 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__B2 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__B2 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__B2 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__C (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__B (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__B2 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__C (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__A1 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__A2 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__A1 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__A1 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__A2 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A1 (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__A3 (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__B (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__A1 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__A1 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__C (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__C (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__B2 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__B2 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__B1 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__B2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A1 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A1 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__B (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A1 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A1 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__A2 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A2 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A2 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A2 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__B1 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__B1 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A1 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A2 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__B (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__B (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__B (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__B (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__B (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__A2 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__C (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__B (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__A1 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__B (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__I (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A1 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__C (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A2 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__B2 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__B2 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__B2 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__B2 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__B2 (.I(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__A2 (.I(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A2 (.I(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__B2 (.I(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__A1 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A1 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A1 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A1 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__B1 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__B1 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__B1 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__B1 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__B2 (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__B1 (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__A2 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__B2 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__B2 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__B2 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__A1 (.I(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__A1 (.I(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__A1 (.I(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__A1 (.I(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A1 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__A2 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__B2 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A2 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__A2 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__B (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A2 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__C (.I(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__A1 (.I(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7751__A1 (.I(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__A1 (.I(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A2 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A2 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A2 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__A2 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__B (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__C (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A2 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__A1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__I (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A2 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A1 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__A2 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A1 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A2 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A2 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A2 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7751__B (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A2 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__A3 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__B2 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__B1 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__B2 (.I(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__B2 (.I(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__B2 (.I(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__B2 (.I(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__B (.I(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__B (.I(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__B (.I(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__B (.I(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A2 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A3 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A2 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__A1 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A1 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A1 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A1 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__A1 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__I (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A2 (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A1 (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__A1 (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7500__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A2 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__A2 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A1 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__B (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__A2 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__B1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__B1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__B2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__B (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A2 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__B (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A3 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A1 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__A1 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A2 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__A2 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__B (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A3 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__A2 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A2 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A2 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__C (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__B (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__B2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__B2 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__B1 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A1 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A1 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A1 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__A1 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__A1 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__A1 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A1 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A1 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__A1 (.I(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__B2 (.I(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A1 (.I(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__A1 (.I(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__A1 (.I(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__A1 (.I(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__A2 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A2 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__B1 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A2 (.I(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__A2 (.I(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__A1 (.I(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__B2 (.I(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__A1 (.I(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__B (.I(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__B1 (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A1 (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__A1 (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__A1 (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__A1 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__A2 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7562__B (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__B2 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__B2 (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__C1 (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__I (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A1 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__A1 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A1 (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A2 (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__A2 (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__A2 (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A2 (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A2 (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__A1 (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__I (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A1 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__C (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A1 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7583__A1 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__C (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__B (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__B (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__B (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__B (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__B (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__B1 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__B (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7610__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__A2 (.I(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__B1 (.I(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__A2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__B2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7652__I (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__A2 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A2 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__A2 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__A2 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A2 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A2 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A2 (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A3 (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A2 (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__B2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__B1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__A1 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A1 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__C (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__B1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A1 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__A1 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A1 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A1 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__A1 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A1 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A3 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A2 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A2 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__B1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__C (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__C (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__C (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__C (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__B (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__C (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__B (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A1 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A1 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__A1 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A1 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__A3 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__B (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__C (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__B (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__B (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__B (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__B (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A1 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__A1 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A1 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__A1 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__B2 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__B1 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__B1 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A1 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__C (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A1 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A1 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__B (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__C (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__B (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__B (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A1 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A1 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__B (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A2 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__B (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__C (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A1 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__A2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__C (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__B (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__A2 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A2 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__A1 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__B1 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__B2 (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__C (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__C (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A1 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A2 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__C (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__C (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__C (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__C (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__B1 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__B2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__B (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__C (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A2 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__A1 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__A1 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A1 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__B (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__A1 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A1 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A1 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__I (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__C (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__B (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__B (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__C (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A1 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__B2 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__B (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__B (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__B (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__B (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__C (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__C (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A1 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__I (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A4 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A3 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A2 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__C (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A4 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A2 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A2 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A2 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A2 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__B (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__I (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A2 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__C (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__I (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__I (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__I (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__A2 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__A2 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A1 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A2 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A2 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A2 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A2 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A2 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__B (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__C (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__C (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__I (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A1 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A1 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A2 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A2 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A1 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A1 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A1 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A1 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__B (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__B1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A2 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__B1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__B2 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__B1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__I (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__A2 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__A2 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__B1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__B (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__B (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__B (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__B (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__C (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__B1 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__B (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__B (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__C (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A2 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__B (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A3 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__A2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A1 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__A1 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A1 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__A1 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__C (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__B2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__B2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__A1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__C (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__B (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A2 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A1 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__B (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__A2 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__B (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__B (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__B (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A2 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__B1 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__C (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__B (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__B (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__C (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__B (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__C (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__C (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__B2 (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__C (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__C (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__C (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__C (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__B (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__B1 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__B (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A1 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__B2 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A2 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__C (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__B (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__B (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__B (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__B (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__B (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__A2 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__A2 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__I (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__I (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__A2 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__A2 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A2 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__A2 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__B (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__A2 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__A2 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__I (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__I (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A2 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A2 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A2 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A2 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__A2 (.I(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__A2 (.I(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__A2 (.I(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__A2 (.I(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__A1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__A1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__A2 (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__A2 (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__A2 (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A2 (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__B (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A2 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A3 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A2 (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8070__A4 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__I (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__I (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__B (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__I (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__I (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__I (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__A1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__A1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8419__B2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__C (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__C (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__C (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__I (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__B (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__B (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__C (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__I (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A1 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__B2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__B (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__B2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__A2 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A2 (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__A1 (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A1 (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A1 (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__A1 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__B2 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__A1 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__I (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__A2 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__A2 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__I (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A2 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__B1 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A2 (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8426__A2 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__A2 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__A2 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__A2 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__I (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__I (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A2 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__A2 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__A2 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__I (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A2 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__A2 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__A2 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A2 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__A1 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A1 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__B2 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A1 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8419__A1 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__A1 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__B2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__A1 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__B2 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__B2 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__B2 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__B2 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__B (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__A2 (.I(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__C (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__A1 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A1 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__C (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__A1 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__B2 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__B2 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A1 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A2 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__B2 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__B2 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__B2 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__I (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__B2 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__B2 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__B2 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__B2 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__C (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__B1 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A2 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__B1 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__B2 (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__A1 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__I (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__I (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__C (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__B (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A1 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A1 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__A2 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__A2 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__A1 (.I(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__A1 (.I(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__A1 (.I(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__A1 (.I(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__A2 (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__A2 (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__C (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__B (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A2 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A2 (.I(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__B1 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__B (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__B1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__B1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A2 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__B1 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A2 (.I(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__A1 (.I(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A3 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__A2 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__A1 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__A3 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__A2 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A3 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8280__B1 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A2 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A3 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__A2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__B1 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__A2 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__B2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__A3 (.I(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__A1 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A1 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A1 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A1 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A2 (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A2 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__A2 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A2 (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__A2 (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__A2 (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__B1 (.I(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__A1 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__A1 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A1 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A1 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__A2 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__I (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A2 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A2 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__B2 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__A2 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A2 (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A2 (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__A2 (.I(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__C (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__C (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A1 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__C (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A2 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8291__A2 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__A2 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A2 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A2 (.I(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__B1 (.I(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__B (.I(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__C (.I(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__C (.I(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__C (.I(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__C (.I(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A1 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A1 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__A2 (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__A1 (.I(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__A2 (.I(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A1 (.I(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__A2 (.I(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__A3 (.I(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A2 (.I(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A2 (.I(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A2 (.I(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__A2 (.I(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__A2 (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__B (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A2 (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__A4 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A2 (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A2 (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__B2 (.I(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__A2 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__A2 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A2 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A2 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A2 (.I(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A2 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A2 (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A2 (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__B2 (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__A2 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__A2 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__A2 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8397__I0 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__B (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__B (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__B (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A1 (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A1 (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A1 (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A1 (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__A2 (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__B (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8397__I1 (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A2 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A2 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__A2 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__A2 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A2 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__B1 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__C (.I(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__B1 (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A2 (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A2 (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__I (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A2 (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__A2 (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A2 (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A2 (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__B1 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8454__A2 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A2 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__A2 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A1 (.I(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__A1 (.I(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__A1 (.I(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A1 (.I(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A2 (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A2 (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A2 (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A2 (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__A1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__B2 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__A1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__A1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__B2 (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A2 (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A2 (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A2 (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A1 (.I(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A2 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A3 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__A1 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A3 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A2 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A4 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__A3 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__B (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__B2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__B (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__B (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__B1 (.I(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__B1 (.I(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__B1 (.I(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A2 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__A1 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A1 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A1 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__B (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__A1 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__A1 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__A2 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A1 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__A1 (.I(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A2 (.I(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A2 (.I(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A3 (.I(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__A2 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__A2 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__A1 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A2 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__C (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__B1 (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A1 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__A2 (.I(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A2 (.I(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__B1 (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__B1 (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__B1 (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__A1 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__A2 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__A2 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__A4 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__B (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A2 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__B2 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A3 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__A3 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__B (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__I (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__A1 (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__A1 (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__A1 (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__A2 (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__C (.I(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__A2 (.I(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__B (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__B (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__I (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__B2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__B2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__B2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__B (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__S0 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__S0 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__S0 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__I (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__S0 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A1 (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A1 (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__S (.I(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__S (.I(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__S (.I(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__I (.I(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__S1 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__I (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__S (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__I (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__S1 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__S (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__I (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A1 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__S1 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A1 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__I (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A1 (.I(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A2 (.I(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__I (.I(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A2 (.I(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__I (.I(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A1 (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__I (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__I (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__I (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A1 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A1 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__I (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__I (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__I (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A1 (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8347__I (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__I (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__I (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A2 (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A2 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__I (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__I (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A2 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A1 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A1 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A3 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__I (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__I (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A1 (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A1 (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A1 (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A2 (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A2 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A1 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__B2 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A2 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A2 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A2 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__B2 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__B2 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A2 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A1 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A2 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__C (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__I (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A1 (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__A1 (.I(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__I (.I(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A1 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A1 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A1 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__I (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__I (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A4 (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A1 (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__A1 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__B2 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__A1 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A2 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__C (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A1 (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A2 (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A2 (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__I (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__I (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A1 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A2 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A1 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__I (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A1 (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A2 (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A2 (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A2 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__I (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A2 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__B (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__I (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A2 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__I (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__I (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A2 (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__I (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A1 (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__I (.I(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A2 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__I (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__I (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A1 (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A1 (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A2 (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__B1 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A2 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__I (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__B2 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A3 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A2 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A2 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A2 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A3 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__I (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__C (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__I (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A1 (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__I (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A2 (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__I (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A1 (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__I (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__I (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A2 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__B2 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A3 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A1 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A2 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__I (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__I (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A2 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A2 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__I (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__I (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__I (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__I (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__I (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A2 (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A1 (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A1 (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__I (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A3 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A3 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A3 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A2 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__I (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A1 (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A3 (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A2 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A3 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A3 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A2 (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__I (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A1 (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A1 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A3 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A2 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A3 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__A1 (.I(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__I (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A1 (.I(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__I (.I(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A1 (.I(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__B2 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A2 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A1 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__I (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A1 (.I(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A1 (.I(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A3 (.I(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A1 (.I(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__I (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A3 (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__I (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A1 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__B2 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A2 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A2 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__I (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__S0 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A2 (.I(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A2 (.I(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__I (.I(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A2 (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A2 (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__I (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__I (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__I (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A3 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__I (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A2 (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__I (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A1 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__I (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A1 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__I (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__I (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A1 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__I (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__A1 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__I (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A2 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A1 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A1 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A1 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A4 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A2 (.I(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A3 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__I (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A3 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__I (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__I (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A1 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__B2 (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A1 (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__B (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A2 (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__I (.I(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__I (.I(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A4 (.I(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__I (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__I (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__I (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__B (.I(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A1 (.I(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A1 (.I(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A1 (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A1 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A1 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A2 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A2 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__C (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__I (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__I (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A2 (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A2 (.I(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A3 (.I(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A3 (.I(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A3 (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__I (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A2 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__A1 (.I(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A2 (.I(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A2 (.I(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A1 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A1 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__I (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__B (.I(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A1 (.I(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__A1 (.I(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A1 (.I(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A1 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__B2 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A2 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__B (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__B (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__I (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__B2 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__I (.I(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__I (.I(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__I (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A1 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__S1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__I (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__S1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__S (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A2 (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A2 (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A2 (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A2 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__B2 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__I (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__I (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__I (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__B1 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A2 (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__B2 (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A2 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__I (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I (.I(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A1 (.I(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__B2 (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__B2 (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__B2 (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A2 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__I (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__A2 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A2 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A1 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A2 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A2 (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__I (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__I (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__I0 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__B (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A2 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__C (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__I (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A2 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A1 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A1 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__I (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A2 (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A2 (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__I (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__I (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__I (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__I (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A1 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A1 (.I(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__I (.I(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__I (.I(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__I (.I(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__B (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__B (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__B (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__B (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__B (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A1 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__I (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A3 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__S1 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__S (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__S1 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__S (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__A2 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A2 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A2 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A1 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__I (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A2 (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A2 (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__I (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A1 (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__B2 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A4 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__I (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__A2 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A2 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A2 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__I (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__I (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A1 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A1 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A1 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__I (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__I (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A2 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A1 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A3 (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A3 (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A1 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A1 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A1 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__I (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A2 (.I(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A2 (.I(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A2 (.I(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__A1 (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A1 (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A2 (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__B (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__B (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__B (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__B1 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__B (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__C (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__B2 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A1 (.I(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A1 (.I(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A1 (.I(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__C (.I(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__B (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__C (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A1 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A2 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A2 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A1 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A1 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__I (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A1 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__A1 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A1 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__B (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__I (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__I (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A3 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__I (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__I (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A4 (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__I (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__I (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__C2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__B2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__B2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__I (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A2 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__A2 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A1 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A1 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__I (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__I (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__B (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A3 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__C (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__C (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__B (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A2 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__I (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A2 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A1 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__B (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A2 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__I (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__B (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A1 (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__A1 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A1 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A1 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A1 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__I (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A1 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A2 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A1 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__I (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__B (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A2 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A1 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__I (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A2 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__B (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__I (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A1 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A2 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__I (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__C (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__I (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__C (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__B (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A1 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__A1 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A2 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A1 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__I (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__I (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A1 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__I (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A1 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A2 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__I (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__I (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A2 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__I (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A1 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A2 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A1 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A3 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__A2 (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A1 (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A3 (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A1 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A1 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A2 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__I (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__I (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__I (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A1 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A1 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__I (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__B2 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A1 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A1 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__I (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A4 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__I (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__I (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__I (.I(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A1 (.I(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A3 (.I(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A2 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A2 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A2 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A2 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A2 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A3 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__I (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__B2 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__I (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A1 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A1 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__B2 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A1 (.I(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A1 (.I(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__B2 (.I(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A2 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A2 (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A2 (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__I (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A2 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A3 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7806__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__I (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A3 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A3 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A1 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__I (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__A1 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A3 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A2 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A3 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__I (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A2 (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__A2 (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__B2 (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A4 (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__B2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__B2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__B2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A2 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__B1 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__A2 (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A2 (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A1 (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A2 (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A2 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__B2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A1 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A2 (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A1 (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A1 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__I (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A2 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__I (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A1 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A1 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A1 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__A2 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A2 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__B2 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__I (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A1 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A1 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__I (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A1 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__I (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__B2 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__I (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A2 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__I (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__I (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A1 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A2 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__I (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__B2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A1 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A1 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A2 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__I (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A2 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A1 (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A4 (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A2 (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__A1 (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A2 (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__I (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__I (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A1 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__B (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A1 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__I (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A1 (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A1 (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A1 (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__I (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A1 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A1 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__I (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__B (.I(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__A2 (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__C (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A1 (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A2 (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A1 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__I (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__B (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__B (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__I (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A1 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__B2 (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A1 (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A1 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A3 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__I (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A1 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A1 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A1 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__B (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A3 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A2 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A2 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__B (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A3 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A3 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A1 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__I (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A2 (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A1 (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__I (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__I (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A2 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A1 (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A1 (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__I (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A1 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__B (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__I (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__I (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__A2 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__I (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A1 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A2 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__I (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__I (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__I (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A3 (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__I (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__I (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__B2 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A3 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__I (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7685__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A2 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__A1 (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__A1 (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__A1 (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__I (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__A1 (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__I (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__I (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__I (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A2 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__I (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A1 (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__A1 (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__I (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__I (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__S (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__S (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__S (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__I (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__I (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__I (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__B (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__I (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__I (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__B2 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__I (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__I (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A1 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__I0 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__I1 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__A1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__I0 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__I1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__I0 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__I1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I0 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__I1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__I0 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__I0 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__I1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__I0 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A1 (.I(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__I0 (.I(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A1 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__I0 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__I1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__I3 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__I1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__I3 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__I1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__I3 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__I3 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__I1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I3 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__I1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__I3 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__I1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__I3 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__B2 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__I2 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__B1 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A1 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__B1 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__A1 (.I(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__B1 (.I(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__A1 (.I(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__B1 (.I(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__B1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__A1 (.I(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__A1 (.I(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A1 (.I(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A2 (.I(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__B1 (.I(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__B1 (.I(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__B1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__B1 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A1 (.I(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A2 (.I(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__B (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__B2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__A3 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8220__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__A3 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8426__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8761__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8758__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8764__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8633__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8635__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8634__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8637__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8639__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8852__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8769__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8853__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8856__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8851__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8850__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8862__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__CLK (.I(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__CLK (.I(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8801__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8802__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__CLK (.I(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__CLK (.I(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__CLK (.I(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__CLK (.I(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8834__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8819__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8694__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8725__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8840__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8833__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8717__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8684__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8674__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8828__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8821__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8820__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8843__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8830__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8726__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8842__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8837__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8813__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8838__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8831__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8829__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8664__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8657__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8816__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8836__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8666__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8704__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8796__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8797__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8874__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8875__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8884__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8882__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8871__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8876__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8724__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8730__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8685__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8845__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8826__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8827__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8825__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8846__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8848__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8719__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8844__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8823__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8822__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8751__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8753__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8737__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8734__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8736__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8879__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8743__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8716__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8870__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8812__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8868__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8867__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8747__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8744__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8863__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8715__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8869__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8864__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8805__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__CLK (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__CLK (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8877__CLK (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8880__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_3_0_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8780__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8766__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8786__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8788__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8854__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__CLK (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_1_wb_clk_i_I (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_opt_1_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_1_wb_clk_i_I (.I(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__CLK (.I(clknet_opt_2_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__CLK (.I(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net88;
 assign io_oeb[13] = net93;
 assign io_oeb[14] = net53;
 assign io_oeb[15] = net54;
 assign io_oeb[16] = net55;
 assign io_oeb[17] = net56;
 assign io_oeb[18] = net57;
 assign io_oeb[19] = net58;
 assign io_oeb[1] = net89;
 assign io_oeb[20] = net59;
 assign io_oeb[21] = net60;
 assign io_oeb[22] = net61;
 assign io_oeb[23] = net62;
 assign io_oeb[24] = net63;
 assign io_oeb[25] = net64;
 assign io_oeb[26] = net65;
 assign io_oeb[27] = net66;
 assign io_oeb[28] = net67;
 assign io_oeb[29] = net68;
 assign io_oeb[2] = net90;
 assign io_oeb[30] = net69;
 assign io_oeb[31] = net70;
 assign io_oeb[32] = net71;
 assign io_oeb[33] = net72;
 assign io_oeb[34] = net73;
 assign io_oeb[35] = net74;
 assign io_oeb[36] = net75;
 assign io_oeb[37] = net76;
 assign io_oeb[3] = net91;
 assign io_oeb[4] = net92;
 assign io_out[0] = net77;
 assign io_out[13] = net82;
 assign io_out[1] = net78;
 assign io_out[2] = net79;
 assign io_out[33] = net83;
 assign io_out[34] = net84;
 assign io_out[35] = net85;
 assign io_out[36] = net86;
 assign io_out[37] = net87;
 assign io_out[3] = net80;
 assign io_out[4] = net81;
endmodule

