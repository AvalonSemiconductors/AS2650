VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO serial_ports
  CLASS BLOCK ;
  FOREIGN serial_ports ;
  ORIGIN 0.000 0.000 ;
  SIZE 275.000 BY 275.000 ;
  PIN RXD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 0.000 193.200 4.000 ;
    END
  END RXD
  PIN TXD
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 0.000 170.800 4.000 ;
    END
  END TXD
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 15.680 275.000 16.240 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 29.120 275.000 29.680 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 42.560 275.000 43.120 ;
    END
  END addr[2]
  PIN bus_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 4.000 ;
    END
  END bus_cyc
  PIN bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 0.000 238.000 4.000 ;
    END
  END bus_we
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 56.000 275.000 56.560 ;
    END
  END data_in[0]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 69.440 275.000 70.000 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 82.880 275.000 83.440 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 96.320 275.000 96.880 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 109.760 275.000 110.320 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 123.200 275.000 123.760 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 136.640 275.000 137.200 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 150.080 275.000 150.640 ;
    END
  END data_in[7]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 163.520 275.000 164.080 ;
    END
  END data_out[0]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 176.960 275.000 177.520 ;
    END
  END data_out[1]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 190.400 275.000 190.960 ;
    END
  END data_out[2]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 203.840 275.000 204.400 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 217.280 275.000 217.840 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 230.720 275.000 231.280 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 244.160 275.000 244.720 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 271.000 257.600 275.000 258.160 ;
    END
  END data_out[7]
  PIN io_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END io_in
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 0.000 103.600 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 0.000 126.000 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 0.000 148.400 4.000 ;
    END
  END io_oeb[2]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 0.000 36.400 4.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END io_out[2]
  PIN irq3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 0.000 260.400 4.000 ;
    END
  END irq3
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 271.000 206.640 275.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 259.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 259.020 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 259.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 259.020 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 271.000 68.880 275.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Pwell ;
        RECT 6.290 256.960 268.670 259.150 ;
      LAYER Nwell ;
        RECT 6.290 252.765 268.670 256.960 ;
        RECT 6.290 252.640 88.305 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 268.670 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 155.720 249.120 ;
        RECT 6.290 244.800 268.670 248.995 ;
      LAYER Pwell ;
        RECT 6.290 241.280 268.670 244.800 ;
      LAYER Nwell ;
        RECT 6.290 237.085 268.670 241.280 ;
        RECT 6.290 236.960 52.465 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 268.670 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 68.705 233.440 ;
        RECT 6.290 229.120 268.670 233.315 ;
      LAYER Pwell ;
        RECT 6.290 225.600 268.670 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 131.985 225.600 ;
        RECT 6.290 221.405 268.670 225.475 ;
        RECT 6.290 221.280 37.905 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 268.670 221.280 ;
      LAYER Nwell ;
        RECT 6.290 213.565 268.670 217.760 ;
        RECT 6.290 213.440 77.665 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 268.670 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 135.345 209.920 ;
        RECT 6.290 205.725 268.670 209.795 ;
        RECT 6.290 205.600 40.705 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 268.670 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 113.830 202.080 ;
        RECT 6.290 197.885 268.670 201.955 ;
        RECT 6.290 197.760 32.305 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 268.670 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 64.225 194.240 ;
        RECT 6.290 190.045 268.670 194.115 ;
        RECT 6.290 189.920 168.945 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 268.670 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 12.705 186.400 ;
        RECT 6.290 182.205 268.670 186.275 ;
        RECT 6.290 182.080 236.705 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 268.670 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 180.705 178.560 ;
        RECT 6.290 174.365 268.670 178.435 ;
        RECT 6.290 174.240 12.705 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 268.670 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 108.465 170.720 ;
        RECT 6.290 166.525 268.670 170.595 ;
        RECT 6.290 166.400 133.880 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 268.670 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 12.705 162.880 ;
        RECT 6.290 158.685 268.670 162.755 ;
        RECT 6.290 158.560 53.025 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 268.670 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 81.350 155.040 ;
        RECT 6.290 150.845 268.670 154.915 ;
        RECT 6.290 150.720 12.705 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 268.670 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 70.945 147.200 ;
        RECT 6.290 143.005 268.670 147.075 ;
        RECT 6.290 142.880 161.105 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 268.670 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 12.705 139.360 ;
        RECT 6.290 135.165 268.670 139.235 ;
        RECT 6.290 135.040 71.505 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 268.670 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 143.960 131.520 ;
        RECT 6.290 127.325 268.670 131.395 ;
        RECT 6.290 127.200 159.985 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 268.670 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 12.705 123.680 ;
        RECT 6.290 119.485 268.670 123.555 ;
        RECT 6.290 119.360 73.745 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 268.670 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 261.000 115.840 ;
        RECT 6.290 111.645 268.670 115.715 ;
        RECT 6.290 111.520 12.705 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 268.670 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 71.505 108.000 ;
        RECT 6.290 103.805 268.670 107.875 ;
        RECT 6.290 103.680 54.145 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 268.670 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 91.105 100.160 ;
        RECT 6.290 95.965 268.670 100.035 ;
        RECT 6.290 95.840 12.705 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 268.670 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 31.275 92.320 ;
        RECT 6.290 88.125 268.670 92.195 ;
        RECT 6.290 88.000 93.345 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 268.670 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 12.705 84.480 ;
        RECT 6.290 80.285 268.670 84.355 ;
        RECT 6.290 80.160 51.905 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 268.670 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 97.825 76.640 ;
        RECT 6.290 72.445 268.670 76.515 ;
        RECT 6.290 72.320 200.070 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 268.670 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 12.705 68.800 ;
        RECT 6.290 64.605 268.670 68.675 ;
        RECT 6.290 64.480 157.745 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 268.670 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 255.745 60.960 ;
        RECT 6.290 56.765 268.670 60.835 ;
        RECT 6.290 56.640 12.705 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 268.670 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 103.985 53.120 ;
        RECT 6.290 48.925 268.670 52.995 ;
        RECT 6.290 48.800 20.200 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 268.670 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 227.280 45.280 ;
        RECT 6.290 41.085 268.670 45.155 ;
        RECT 6.290 40.960 40.705 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 268.670 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 30.625 37.440 ;
        RECT 6.290 33.245 268.670 37.315 ;
        RECT 6.290 33.120 71.505 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 268.670 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 173.985 29.600 ;
        RECT 6.290 25.405 268.670 29.475 ;
        RECT 6.290 25.280 49.105 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 268.670 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 103.985 21.760 ;
        RECT 6.290 17.565 268.670 21.635 ;
        RECT 6.290 17.440 126.945 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 268.670 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 268.240 259.020 ;
      LAYER Metal2 ;
        RECT 8.540 270.700 68.020 271.000 ;
        RECT 69.180 270.700 205.780 271.000 ;
        RECT 206.940 270.700 266.980 271.000 ;
        RECT 8.540 4.300 266.980 270.700 ;
        RECT 8.540 4.000 13.140 4.300 ;
        RECT 14.300 4.000 35.540 4.300 ;
        RECT 36.700 4.000 57.940 4.300 ;
        RECT 59.100 4.000 80.340 4.300 ;
        RECT 81.500 4.000 102.740 4.300 ;
        RECT 103.900 4.000 125.140 4.300 ;
        RECT 126.300 4.000 147.540 4.300 ;
        RECT 148.700 4.000 169.940 4.300 ;
        RECT 171.100 4.000 192.340 4.300 ;
        RECT 193.500 4.000 214.740 4.300 ;
        RECT 215.900 4.000 237.140 4.300 ;
        RECT 238.300 4.000 259.540 4.300 ;
        RECT 260.700 4.000 266.980 4.300 ;
      LAYER Metal3 ;
        RECT 8.490 258.460 271.000 258.860 ;
        RECT 8.490 257.300 270.700 258.460 ;
        RECT 8.490 245.020 271.000 257.300 ;
        RECT 8.490 243.860 270.700 245.020 ;
        RECT 8.490 231.580 271.000 243.860 ;
        RECT 8.490 230.420 270.700 231.580 ;
        RECT 8.490 218.140 271.000 230.420 ;
        RECT 8.490 216.980 270.700 218.140 ;
        RECT 8.490 204.700 271.000 216.980 ;
        RECT 8.490 203.540 270.700 204.700 ;
        RECT 8.490 191.260 271.000 203.540 ;
        RECT 8.490 190.100 270.700 191.260 ;
        RECT 8.490 177.820 271.000 190.100 ;
        RECT 8.490 176.660 270.700 177.820 ;
        RECT 8.490 164.380 271.000 176.660 ;
        RECT 8.490 163.220 270.700 164.380 ;
        RECT 8.490 150.940 271.000 163.220 ;
        RECT 8.490 149.780 270.700 150.940 ;
        RECT 8.490 137.500 271.000 149.780 ;
        RECT 8.490 136.340 270.700 137.500 ;
        RECT 8.490 124.060 271.000 136.340 ;
        RECT 8.490 122.900 270.700 124.060 ;
        RECT 8.490 110.620 271.000 122.900 ;
        RECT 8.490 109.460 270.700 110.620 ;
        RECT 8.490 97.180 271.000 109.460 ;
        RECT 8.490 96.020 270.700 97.180 ;
        RECT 8.490 83.740 271.000 96.020 ;
        RECT 8.490 82.580 270.700 83.740 ;
        RECT 8.490 70.300 271.000 82.580 ;
        RECT 8.490 69.140 270.700 70.300 ;
        RECT 8.490 56.860 271.000 69.140 ;
        RECT 8.490 55.700 270.700 56.860 ;
        RECT 8.490 43.420 271.000 55.700 ;
        RECT 8.490 42.260 270.700 43.420 ;
        RECT 8.490 29.980 271.000 42.260 ;
        RECT 8.490 28.820 270.700 29.980 ;
        RECT 8.490 16.540 271.000 28.820 ;
        RECT 8.490 15.540 270.700 16.540 ;
      LAYER Metal4 ;
        RECT 109.340 16.890 175.540 252.470 ;
        RECT 177.740 16.890 232.260 252.470 ;
  END
END serial_ports
END LIBRARY

