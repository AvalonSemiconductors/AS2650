* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i wb_rst_i
XFILLER_79_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6209__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7406__A1 _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7957__A2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7963_ _1378_ _2173_ _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5968__A1 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6914_ _2350_ _2351_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7894_ as2650.stack\[4\]\[14\] _1266_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8657__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6845_ _2085_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8382__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7684__C _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6776_ _1400_ _2082_ _2219_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8515_ _1297_ _0462_ _3816_ _3832_ _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5727_ _1249_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8446_ _1388_ _1391_ _1616_ _3775_ _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5658_ _1211_ _1169_ _1214_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4609_ _4171_ _4091_ _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8377_ _2068_ _3701_ _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _4158_ _1156_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7328_ _2743_ _2710_ _2744_ _2745_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7645__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7645__B2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7259_ _2638_ _2678_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7948__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6620__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6384__A1 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7166__I _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8125__A2 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6136__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6687__A2 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7636__A1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7636__B2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5414__I _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__C _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8061__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6611__A2 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4960_ _4162_ _0511_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7785__B _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _0485_ _0412_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _3954_ _2091_ _2092_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5178__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6561_ _2031_ _1652_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_125_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8116__A2 _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8300_ _3642_ _3643_ _2131_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5512_ as2650.stack\[0\]\[2\] _1090_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6127__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6492_ _1970_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8231_ _3900_ _3577_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ _3880_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__I0 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8162_ _2824_ _3510_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5374_ as2650.r123\[0\]\[4\] _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7113_ _1014_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7627__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4325_ _3904_ _3905_ _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8093_ net31 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7044_ _2460_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6850__A2 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4861__A1 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8052__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8052__B2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7946_ as2650.stack\[7\]\[5\] _3300_ _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7877_ _1199_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5994__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6828_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8303__C _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _0457_ _2194_ _2206_ _2207_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4916__A2 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8107__A2 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6118__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6669__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5943__B _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8429_ _1495_ _2337_ _3759_ _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7714__I _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5877__B1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7094__A2 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4852__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8043__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6054__B1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6065__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5580__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7306__B1 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__A1 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7609__B2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5883__A3 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7085__A2 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8282__A1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5090_ _0687_ _0601_ _0587_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5096__A1 _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8034__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7800_ _0413_ _3201_ _1494_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8780_ _0257_ clknet_leaf_28_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5992_ _1509_ _0618_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7731_ _1379_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4943_ _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8337__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7662_ _2139_ _2385_ _2443_ _3067_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6348__A1 _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4874_ _0294_ _4156_ _4256_ _0289_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6613_ as2650.cycle\[7\] _3929_ _2072_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6899__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7593_ _3003_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6544_ _0584_ _1656_ _2008_ as2650.r123_2\[1\]\[4\] _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7848__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6475_ _1837_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8214_ _2911_ _3560_ _2912_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5426_ _0889_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8145_ _3336_ _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5357_ _4136_ _0857_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ as2650.cycle\[7\] _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8273__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7076__A2 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8076_ _3330_ _3414_ _3427_ _2226_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5288_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5087__A1 _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5989__I _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7027_ _1634_ _2269_ _1410_ _1421_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_112_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A1 _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6587__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7929_ _3285_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7709__I _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7000__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5562__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8500__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6511__A1 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6814__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8208__C _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8016__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4308__I as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6578__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7782__C _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6750__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5553__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4590_ _3918_ _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6260_ _4212_ _0740_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6502__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5856__A3 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6191_ _3875_ _4206_ _1665_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8255__A1 _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5142_ as2650.r123\[0\]\[6\] as2650.r123_2\[0\]\[6\] _3851_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5069__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5073_ _0652_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6569__A1 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7230__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5975_ _3924_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8763_ _0240_ clknet_leaf_35_wb_clk_i as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5241__A1 _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5241__B2 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7714_ _3120_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8694_ _0171_ clknet_leaf_0_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4857_ _3909_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7645_ _2137_ _2437_ _2444_ _3053_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7576_ _0948_ _2529_ _2968_ _2527_ _2987_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4788_ _0379_ _0382_ _0385_ _0377_ _0388_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6527_ _3849_ _2005_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7264__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6458_ _0646_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5409_ _0998_ _0866_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6389_ _1850_ _1852_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_47_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8246__A1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7049__A2 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8128_ _3448_ _3476_ _3449_ _3477_ _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5940__C _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4837__B _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8059_ _2644_ _3381_ _2690_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6608__I _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8261__A4 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7757__B1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7221__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4586__A3 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6732__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5535__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4338__A3 _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6499__B _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7174__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7288__A2 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8237__A1 _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__I _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6799__A1 _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5223__A1 _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5760_ as2650.stack\[4\]\[7\] _1277_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4711_ _4005_ _4083_ _4086_ _4089_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_72_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7793__B _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ as2650.stack\[2\]\[1\] _1195_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7430_ _2845_ _2799_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4642_ _4221_ _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _2730_ _0543_ _2777_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4734__B1 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4573_ _4136_ _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6312_ _1793_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8476__A1 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7292_ _2377_ _2710_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6243_ _1728_ _1729_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8228__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ _4057_ _1660_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5125_ _0710_ _4060_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7451__A2 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5056_ _0370_ _0563_ _0571_ _0654_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5462__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7687__C _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8400__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5214__A1 _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8746_ _0223_ clknet_leaf_42_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6962__A1 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5958_ _1456_ _0544_ _0690_ _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6962__B2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4909_ _0492_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5889_ _1307_ _1405_ _1406_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8677_ _0154_ clknet_leaf_77_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7628_ _1177_ _3012_ _1184_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7559_ _1166_ _2922_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6190__A2 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5507__I _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8467__A1 _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5376__S1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7722__I _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8563__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5205__B2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4803__I1 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4522__S _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8458__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8458__B2 _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6957__B _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7681__A2 _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7433__A2 _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6930_ _2136_ _1482_ _1345_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__A3 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _2303_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7197__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8600_ _0077_ clknet_leaf_34_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5812_ _1310_ _1321_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6792_ _2108_ _2141_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5747__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8531_ _0008_ clknet_leaf_65_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5743_ as2650.stack\[4\]\[0\] _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ _1222_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8462_ _3767_ _3786_ _3791_ _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_124_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7413_ _2827_ _2828_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4625_ _3886_ _4204_ _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8393_ _4097_ _0460_ _3120_ _1530_ _2180_ _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_117_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8449__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7344_ _2716_ as2650.stack\[5\]\[4\] as2650.stack\[4\]\[4\] _2758_ _2762_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4556_ _3964_ _3966_ _3978_ _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6867__B _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8586__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7275_ _1312_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4487_ _4067_ _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7121__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6226_ _1712_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7672__A2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6157_ _1647_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7424__A2 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6227__A3 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ _1162_ _1592_ _1595_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5997__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5435__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _0613_ _4061_ _4115_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7210__C _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__A4 _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7188__A1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5738__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6935__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4946__B1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8729_ _0206_ clknet_leaf_51_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6702__A4 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput20 net20 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput31 net31 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A2 _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8283__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5700__I _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8391__A3 _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7351__A1 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4410_ _3865_ _3939_ _3990_ _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5390_ _0897_ as2650.stack\[1\]\[13\] as2650.stack\[0\]\[13\] _0901_ _0981_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5901__A2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4341_ as2650.ins_reg\[5\] _3921_ _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7103__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8446__A4 _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7060_ _2322_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4272_ _3852_ _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7654__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6011_ _1527_ _1455_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7406__A2 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7962_ _3316_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5610__I _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5968__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6090__A1 as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7030__C _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _1518_ _1606_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7893_ _3260_ _1269_ _3271_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6844_ _1605_ _2286_ _1294_ _2031_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6775_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7590__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8514_ _3212_ _3834_ _3836_ _3833_ _2372_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_91_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5726_ _1237_ _1250_ _1257_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7981__B _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8445_ _1364_ _2085_ _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5657_ as2650.stack\[1\]\[9\] _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7342__B2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _4180_ _4182_ _4183_ _4187_ _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8376_ _3699_ _3710_ _3711_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5588_ _1159_ _1156_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7893__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7327_ _0541_ _0406_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4539_ _3975_ as2650.idx_ctrl\[0\] _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_137_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7645__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7258_ _2573_ _2648_ _2574_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _4050_ _1673_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7189_ _2606_ _2609_ _1323_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8601__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__A3 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__A1 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8751__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6136__A2 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7884__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4698__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7182__I _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7115__C _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7636__A2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5430__I as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4890_ _0426_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7785__C _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7572__A1 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7572__B2 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6560_ _0458_ _0851_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5511_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6491_ _1926_ _1962_ _1971_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6127__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7324__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5442_ _1024_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8230_ _0806_ _0821_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7875__A2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6922__I1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__A1 _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8161_ _2828_ _3442_ _2829_ _2825_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5373_ _0954_ _0934_ _0965_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4324_ _3877_ _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_99_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7112_ _0875_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8092_ _2465_ _3442_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7627__A2 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7043_ _2470_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8624__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4861__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8052__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7945_ _1239_ _3298_ _3303_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8774__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7876_ _3260_ _1578_ _3261_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7012__B1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6827_ _1362_ _2074_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6171__I _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ as2650.r123\[2\]\[3\] _2202_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5709_ _1244_ _1240_ _1245_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6118__A2 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7315__A1 as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6689_ _2074_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8428_ _3729_ _2336_ _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7866__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5877__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5877__B2 _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8359_ net44 _3688_ _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4852__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6054__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6054__B2 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6357__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A1 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A1 _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6109__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7306__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5425__I _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8647__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7609__A2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8282__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8797__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8034__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7793__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7730_ _3131_ _4195_ _3132_ _3135_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4942_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8404__C _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8337__A3 _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7661_ _2662_ _2836_ _3068_ _2885_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7545__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6348__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4873_ _0470_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7545__B2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6612_ _3890_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7592_ as2650.pc\[11\] _1483_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6899__A3 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6543_ _1871_ _2011_ _2018_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7848__A2 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ _1926_ _1955_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8213_ _3510_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5425_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6520__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8144_ _3132_ _2333_ _3490_ _3493_ _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5356_ _0949_ _0866_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6875__B _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8793__D _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4307_ _3887_ _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8273__A2 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8075_ _3420_ _3426_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ as2650.psu\[0\] _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6284__A1 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5087__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7026_ _2451_ _2454_ _2273_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7481__B1 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4834__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6587__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7784__A1 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7928_ _3258_ _3292_ _3293_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7536__A1 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7859_ as2650.stack\[5\]\[8\] _1586_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4414__I _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7725__I _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7839__A2 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6511__A2 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7460__I _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_39_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6814__A3 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8016__A2 _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7775__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7527__A1 _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5002__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6750__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6502__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6190_ _4065_ _1671_ _1675_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _0658_ _0662_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8466__I _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A2 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5072_ _0655_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7303__C _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4816__A2 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5104__B _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8007__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__A2 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6714__I _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8762_ _0239_ clknet_leaf_35_wb_clk_i as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5974_ _1478_ _1481_ _1491_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7713_ _3919_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4925_ as2650.r123\[0\]\[5\] as2650.r123_2\[0\]\[5\] _0365_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7518__A1 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8693_ _0170_ clknet_leaf_80_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7518__B2 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7644_ _1191_ _3052_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4856_ _0425_ _0456_ _4250_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8191__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7575_ _1636_ _2984_ _2986_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4787_ _4121_ _0386_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_105_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6526_ _2004_ _1702_ _1703_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_118_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6457_ _1806_ _1909_ _1911_ _1939_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8494__A2 _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ _0710_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6388_ as2650.r123_2\[2\]\[3\] _1717_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8127_ _0542_ _0556_ _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8246__A2 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5339_ _0859_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6257__A1 _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6257__B2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7454__B1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8058_ _2409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7213__C _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _1037_ _1028_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6009__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7757__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7757__B2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8044__C _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7509__A1 _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4991__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8182__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6732__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6499__C _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4743__A1 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6496__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6799__A2 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__A2 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _0311_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7793__C _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8173__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5690_ _1088_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _4220_ _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4734__A1 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7360_ _2686_ _2734_ _2735_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4572_ _4054_ _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6311_ _1795_ _1796_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7291_ _2707_ _2659_ _2708_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8476__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6242_ _0780_ _0792_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6709__I _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8228__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6173_ _0458_ _1659_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6239__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5124_ _4094_ _0539_ _0720_ _0721_ _4059_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7987__A1 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5055_ _0653_ _0572_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_84_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7451__A3 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5462__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7739__A1 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8400__A2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5214__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8745_ _0222_ clknet_leaf_41_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _1471_ _1472_ _1473_ _1474_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5765__A3 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4973__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4908_ _4022_ _0498_ _0502_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8676_ _0153_ clknet_leaf_2_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5888_ _1007_ _1283_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4899__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7627_ as2650.pc\[12\] _2993_ _3012_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4839_ _4189_ _4177_ _0340_ _4172_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7275__I _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4725__A1 _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _2128_ _2969_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _1955_ _1962_ _1973_ _1988_ _1004_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_101_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7489_ _1158_ _2902_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7978__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6650__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4964__A1 _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4716__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8458__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7913__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_54_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7134__B _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5433__I _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7969__A1 _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__C _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6641__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _2302_ _1296_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7197__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8394__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5811_ _1323_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6791_ _3930_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8530_ _0007_ clknet_leaf_71_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5742_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8146__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8461_ _3788_ _3790_ _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5673_ as2650.r123_2\[3\]\[2\] _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5608__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7412_ as2650.pc\[5\] net1 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4624_ _3913_ _3869_ _3916_ _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8392_ _2182_ _1417_ _2287_ _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5380__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7343_ _2757_ _2759_ _2760_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8449__A2 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4555_ _4131_ _4135_ _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5544__S _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7274_ _2567_ _2692_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _4005_ _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6225_ _1324_ _1711_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7672__A3 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5343__I _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7979__B _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6156_ as2650.r123\[3\]\[4\] _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5107_ _4122_ _0634_ _0700_ _4121_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_44_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6227__A4 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6087_ as2650.stack\[6\]\[8\] _1594_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6632__A1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5435__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _4112_ _0614_ _0624_ _0636_ _4062_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ _1317_ _2411_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5738__A3 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6935__A2 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6902__I _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__A1 _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8728_ _0205_ clknet_leaf_51_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8137__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8659_ _0136_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__I _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6699__A1 _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8530__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5371__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput21 net21 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput43 net43 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5253__I _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8680__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6623__A1 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6084__I _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8376__A1 _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6926__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4332__I as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7351__A2 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5901__A3 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4340_ as2650.ins_reg\[4\] _3868_ as2650.ins_reg\[7\] _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7103__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4271_ _3851_ _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_99_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5665__A2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _1434_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7961_ _3315_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6090__A2 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6912_ _0949_ _2147_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7892_ as2650.stack\[4\]\[13\] _1266_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__A3 _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6843_ _2037_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6722__I _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _3953_ _1405_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7590__A2 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8513_ _0998_ _2367_ _3835_ _1506_ _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ as2650.stack\[3\]\[3\] _1254_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8553__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5338__I as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8444_ _2179_ _1318_ _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5656_ _1134_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5353__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4607_ _4184_ _4185_ _4186_ _4013_ _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8375_ net20 _3704_ _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5587_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7553__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7326_ net9 _0406_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4538_ _4118_ _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6169__I _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7257_ _2636_ _2638_ _2676_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4469_ _4048_ _4049_ _3900_ _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_85_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6853__A1 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ _1657_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7188_ _2215_ _2607_ _2608_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _0840_ _1636_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6605__A1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8070__A3 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6118__B _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6081__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6620__A4 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8358__A1 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__A2 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__B2 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7333__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6788__B _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7097__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6844__A1 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5647__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8061__A3 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8349__A1 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8576__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__A1 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5510_ _1093_ _1085_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6490_ _1959_ _1961_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8521__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ _1025_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8160_ _2812_ _3502_ _3508_ _2595_ _3126_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5886__A2 _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5372_ _0955_ _0936_ _0869_ _0964_ _0861_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_47_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7088__A1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7111_ _2530_ _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4323_ _3876_ _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8091_ _2733_ _3440_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7627__A3 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5638__A2 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7042_ _2469_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6717__I _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5621__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8137__C _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6063__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7260__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7944_ as2650.stack\[7\]\[4\] _3300_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7976__C _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7875_ as2650.stack\[5\]\[13\] _1575_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7012__A1 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ net26 _2269_ _2144_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7563__A2 _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6757_ _2199_ _1895_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ as2650.stack\[2\]\[6\] _1229_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6688_ _0808_ _2123_ _2143_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7315__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8512__A1 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8427_ _1622_ _3718_ _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_137_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5639_ _1202_ _1162_ _1203_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4700__I _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5877__A2 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8358_ _3684_ _0303_ _3696_ _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7309_ _2685_ _2697_ _2726_ _2727_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8289_ _2979_ _3633_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6826__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__I as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8047__C _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8599__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7251__B2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A2 _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5565__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4368__A2 _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7306__A2 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7193__I _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6817__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__A2 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _0543_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7793__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5597__B _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4941_ net9 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__I _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7660_ as2650.pc\[14\] _3055_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ _4196_ _0369_ _0472_ _4000_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7545__A2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6611_ _1314_ _2073_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7591_ _2999_ _3000_ _3001_ _2417_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5020__A3 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6542_ as2650.r123_2\[1\]\[3\] _2015_ _2017_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_9_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6473_ _1954_ _1930_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5616__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8212_ _3407_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5424_ _1009_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8143_ _2493_ _3492_ _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5355_ _0290_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6875__C _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6808__A1 _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4306_ _3886_ _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8074_ _3357_ _3424_ _3425_ _2401_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5286_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7025_ _2452_ _2453_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7481__A1 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6284__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8741__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7481__B2 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6891__B _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7233__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7927_ as2650.stack\[7\]\[12\] _3288_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4598__A2 _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7858_ _1577_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _3908_ _1404_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5547__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7789_ _3181_ _3191_ _3099_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__I _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7472__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5235__B1 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7775__A2 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4589__A2 _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__I _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6820__I _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8614__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__I _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8764__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5140_ _0735_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7463__A1 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6266__A2 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5071_ _0656_ _0663_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8761_ _0238_ clknet_leaf_49_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5973_ _1482_ _1351_ _1486_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_64_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__I _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7712_ _1530_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4924_ as2650.r123\[1\]\[5\] as2650.r123_2\[1\]\[5\] _3855_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8692_ _0169_ clknet_leaf_80_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7643_ _1184_ _1177_ _2994_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8191__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7574_ _2565_ _2968_ _2985_ _2426_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4786_ _0310_ _0314_ _0381_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7047__B _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6525_ _1657_ _1689_ _1705_ _2003_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_88_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _1912_ _1938_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6886__B _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5407_ _0937_ _0992_ _0994_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6387_ _1859_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8126_ _0541_ _0556_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5338_ as2650.r123\[0\]\[2\] _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7454__A1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8057_ _3318_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5269_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7008_ _2309_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7206__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6905__I _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__C _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7757__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__A1 _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6126__B _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__I _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4991__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8182__A2 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6640__I _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6732__A3 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8787__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__A2 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5940__A1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7445__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8516__B as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5759__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6420__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8173__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4640_ _4215_ _4217_ _4219_ _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7920__A2 _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4571_ as2650.r123\[1\]\[0\] _4151_ _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5931__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__A2 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6310_ _0408_ _0526_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7290_ _2707_ _2659_ _2708_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_128_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ _0746_ _0750_ _0791_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6172_ _3967_ _1651_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6239__A2 _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ _4077_ _4109_ _4093_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5054_ _0470_ _0571_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4954__B _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7739__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6947__B1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8744_ _0221_ clknet_leaf_43_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5956_ _0593_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4907_ _0503_ _0505_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8675_ _0152_ clknet_leaf_74_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5887_ _1007_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8164__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7626_ _2134_ _3000_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4838_ _0432_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7372__B1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7911__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7557_ _2552_ _2955_ _2920_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4725__A2 _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4769_ _0289_ _4157_ _4257_ _4196_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ _1922_ _1972_ _1957_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7488_ _1129_ _2866_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7675__A1 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6478__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6439_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5804__I _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4489__A1 _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5150__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8109_ _2133_ _3454_ _3459_ _2485_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7978__A2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7240__B _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4803__I3 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7466__I _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8155__A2 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6166__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7902__A2 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5913__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7666__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__I _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_23_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7969__A2 _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8802__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7150__B _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6641__A2 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4652__A1 _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _1324_ _1328_ _1291_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6790_ _1362_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5741_ _1265_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8146__A2 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8460_ _1018_ _0942_ _3789_ _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5672_ _1221_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7411_ _1106_ net9 _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ _4202_ _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8391_ _1375_ _3720_ _3722_ _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5904__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7342_ _2534_ as2650.stack\[3\]\[4\] as2650.stack\[2\]\[4\] _2668_ _1021_ _2760_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_89_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _4134_ _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8449__A3 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4949__B _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7273_ _2688_ _2691_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_85_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4485_ _3949_ _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5624__I as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8000__I _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6224_ _1702_ _1703_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6155_ _1646_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4891__A1 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8082__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _0555_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6632__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5037_ _4078_ _0635_ _4095_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7188__A3 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6988_ _1617_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8727_ _0204_ clknet_3_0_0_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5939_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8137__A2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4703__I _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8658_ _0135_ clknet_leaf_69_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7345__B1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6699__A2 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7609_ _2053_ _2875_ _2996_ _2620_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8589_ _0066_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5371__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7235__B _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput11 net11 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_108_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5534__I _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput33 net52 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput44 net44 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6320__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5123__A2 _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4882__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8073__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6623__A2 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__A1 _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8376__A2 _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6387__A1 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7887__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6934__I0 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7639__A1 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5444__I _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ as2650.psl\[4\] _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4873__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8064__A1 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6275__I _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7960_ _3308_ _3312_ _3314_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_54_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6911_ _2349_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7891_ _3258_ _1269_ _3270_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8367__A2 _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6842_ _2230_ _2284_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6378__A1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6773_ _1348_ _2214_ _2215_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5050__A1 _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5724_ _1234_ _1250_ _1256_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8512_ _3102_ _3795_ _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8443_ _2302_ _1605_ _3770_ _3772_ _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5655_ _1211_ _1162_ _1212_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4606_ _4171_ _4184_ _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8374_ _3700_ _0805_ _3709_ _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5586_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7055__B _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7325_ _0393_ _0296_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4537_ _3865_ _4050_ _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5105__A2 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7256_ _2648_ _2666_ _2674_ _2675_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_116_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4468_ _3899_ _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ _1688_ _1693_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6853__A2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7187_ _1515_ _2309_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4399_ as2650.ins_reg\[2\] as2650.ins_reg\[3\] _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4864__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6138_ _1617_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7802__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _1097_ _1576_ _1582_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7802__B2 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6118__C _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8358__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5041__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5592__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6916__I0 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7744__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6541__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8294__A1 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8294__B2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6844__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8046__A1 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5280__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6823__I _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7021__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6780__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8521__A2 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5440_ _1026_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6532__A1 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5371_ _0867_ _0961_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5886__A3 _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7110_ _0899_ as2650.stack\[1\]\[0\] as2650.stack\[0\]\[0\] _2531_ _2532_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7088__A2 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4322_ _3874_ _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8090_ _2733_ _3440_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5099__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7041_ _2097_ _2172_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4697__I1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8037__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7322__C _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4518__I _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6934__S _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6599__A1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__A2 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7943_ _1237_ _3298_ _3302_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8434__B _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7874_ _1193_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7012__A2 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6825_ _4204_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5023__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5349__I _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6756_ _0364_ _2194_ _2204_ _2205_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5574__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ _1126_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6687_ _2142_ _2119_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8512__A2 _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8426_ _3738_ _3740_ _3755_ _3756_ _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5638_ as2650.stack\[0\]\[8\] _1121_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ as2650.stack\[1\]\[4\] _1140_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5084__I _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8357_ _1101_ _3685_ _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7079__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8276__A1 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7308_ _2470_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8288_ _2473_ _3630_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6826__A2 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7239_ _2656_ _2658_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7787__B1 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8200__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__I _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6762__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__A2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6514__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8519__B _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6817__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7423__B _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8019__A1 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8019__B2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8543__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5878__B _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7590_ _2389_ _2996_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6753__A1 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ _0482_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5020__A4 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6502__B _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6472_ _1928_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8211_ _3408_ _3556_ _3558_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5423_ _0900_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8258__A1 _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8142_ _2776_ _3491_ _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5354_ _0937_ _0940_ _0945_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4305_ as2650.ins_reg\[4\] _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6808__A2 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8073_ _0397_ _3083_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5285_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4819__A1 _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8148__C _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7024_ _1318_ _2160_ _2438_ _2439_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_64_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7052__C _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7481__A2 _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__A2 as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5492__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6891__C _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8430__A1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7926_ _3283_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7857_ _1161_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6808_ _3932_ _2183_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6744__A1 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5547__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7788_ _0547_ _2214_ _3187_ _3188_ _3190_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _3882_ _2189_ _2190_ _2191_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8409_ _3739_ _1976_ _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8566__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6638__I _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5542__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5235__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5235__B2 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6735__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5717__I _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8488__A1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7160__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7153__B _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5070_ _0664_ _0667_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_69_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8412__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5226__A1 _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6423__B1 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8760_ _0237_ clknet_leaf_43_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6974__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ _1361_ _1489_ _3848_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7711_ _3112_ _3115_ _3117_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4923_ _3845_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8691_ _0168_ clknet_leaf_0_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7642_ _2137_ _3050_ _3000_ _2134_ _2852_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ _0426_ _0432_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8431__C _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7328__B _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7573_ _2567_ _2978_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4785_ _0326_ _0313_ _0380_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4531__I _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ _1812_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8589__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _1915_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5406_ _0882_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6386_ _0456_ _1758_ _1869_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8125_ net52 _3474_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5337_ _0849_ _3991_ _4252_ _0931_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6458__I _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5362__I _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8056_ _3407_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7454__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5268_ _3968_ _3974_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5465__A1 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7007_ _2385_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _0765_ _0767_ _0795_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8403__A1 _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__A1 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__I _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__I _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__A2 _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6126__C _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7909_ _3260_ _1252_ _3280_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__B1 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__I _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7390__A1 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7390__B2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5940__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7142__A1 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7199__I _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4616__I _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6956__A1 _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5759__A2 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__A1 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8173__A3 _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7381__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8731__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4351__I _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4570_ _4150_ _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5931__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7133__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6240_ _0778_ _0779_ _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7684__A2 _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6171_ _1657_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _0714_ _4227_ _0719_ _4210_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5447__A1 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5053_ _0574_ _0576_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8493__I _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4954__C _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6947__A1 _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6947__B2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8743_ _0220_ clknet_leaf_48_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5955_ _0413_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _0503_ _0505_ _4180_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8674_ _0151_ clknet_3_3_0_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5886_ _3867_ _3861_ _3972_ _3918_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_139_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7625_ _3031_ _3034_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4837_ _0342_ _0345_ _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4261__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7556_ _2965_ _2967_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4768_ _4053_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4725__A3 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6897__B _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6507_ _1859_ _1975_ _1986_ _1713_ _1987_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4699_ _0295_ _0297_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7487_ _2865_ _2901_ _2433_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7675__A2 _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6438_ _0626_ _1197_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4489__A2 _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5092__I _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ _1778_ _1803_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8108_ _3454_ _3458_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7427__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__C _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8039_ _1513_ _4244_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4661__A2 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6938__A1 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8754__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7363__A1 _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6166__A2 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8312__B1 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7115__B2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7666__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5216__B _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5730__I _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4346__I as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_63_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4652__A2 _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5601__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7657__I as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__A2 _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _1266_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ as2650.r123_2\[3\]\[1\] _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7354__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7410_ _2777_ _2776_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4622_ _4069_ _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8390_ _3078_ _3721_ _1403_ _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4707__A3 _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7341_ _2716_ as2650.stack\[1\]\[4\] as2650.stack\[0\]\[4\] _2758_ _2759_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4553_ _3968_ _3973_ _4133_ _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7106__A1 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7392__I _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8303__B1 _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7272_ _2642_ _2644_ _2690_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4484_ _4064_ _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5668__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6223_ _1704_ _1706_ _1674_ _1709_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8627__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7409__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ as2650.r123\[3\]\[3\] _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4891__A2 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _0701_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8082__A2 _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6085_ _1590_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5640__I _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6093__A1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6632__A3 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8777__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6672__S _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6987_ _2288_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8726_ _0203_ clknet_leaf_9_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5938_ _0825_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8657_ _0134_ clknet_leaf_69_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5869_ _4076_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7345__B2 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7608_ _3002_ _3016_ _3018_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6699__A3 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8588_ _0065_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8398__I _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7539_ as2650.pc\[9\] _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput12 net12 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput23 net23 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput45 net45 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6320__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8073__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__I _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__A2 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__A1 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6387__A2 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7584__A1 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7336__A1 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7887__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6934__I1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6330__B _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5460__I _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8064__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5822__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4625__A2 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6910_ _4171_ _2348_ _2342_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7890_ as2650.stack\[4\]\[12\] _3266_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6841_ _2232_ _2283_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6378__A2 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7575__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ _2171_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5050__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8511_ _1639_ _2360_ _3833_ _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5723_ as2650.stack\[3\]\[2\] _1254_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8442_ _1311_ _1049_ _2546_ _2599_ _3771_ _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_104_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5654_ as2650.stack\[1\]\[8\] _1146_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7878__A2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4605_ _4166_ _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8373_ _1125_ _3701_ _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5585_ as2650.pc\[8\] _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6550__A2 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4561__A1 _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7324_ _1108_ _2741_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4536_ _4040_ _4047_ _4052_ _4116_ _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_89_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _2186_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _3888_ _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6302__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6894__C _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4313__A1 as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6206_ _4047_ _1690_ _1692_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7186_ _2125_ _2473_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4398_ _3957_ _3964_ _3966_ _3978_ _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_86_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4864__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6137_ _0308_ _1632_ _1635_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__A2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ as2650.stack\[5\]\[2\] _1580_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7297__I _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__I _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5041__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8709_ _0186_ clknet_leaf_38_wb_clk_i as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7869__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6916__I1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7246__B _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5545__I _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6541__A2 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4552__A1 _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7097__A3 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8294__A2 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7760__I _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4304__A1 _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6844__A3 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6376__I _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8046__A2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4607__A2 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7201__S _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5280__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7557__A1 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6044__C _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7309__A1 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7309__B2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6532__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5455__I _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5370_ _0962_ _0917_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5886__A4 _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4321_ _3871_ _3885_ _3901_ _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8285__A2 _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6296__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7040_ _2460_ _2463_ _2467_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8037__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__A1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6599__A2 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7796__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ as2650.stack\[7\]\[3\] _3300_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7548__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7873_ _3258_ _1578_ _3259_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4534__I _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6824_ _3941_ _2149_ _2266_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6755_ as2650.r123\[2\]\[2\] _2202_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4782__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5706_ _1242_ _1240_ _1243_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ _2141_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8425_ _1428_ _3737_ _2267_ _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5637_ _1077_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7720__A1 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8356_ _3682_ _3694_ _3695_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5568_ _1135_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7307_ _2695_ _2715_ _2725_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7079__A3 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4519_ _4099_ _3861_ _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8287_ _3625_ _3627_ _3167_ _3631_ _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7580__I _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5499_ _4081_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7238_ _2558_ _2601_ _2657_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6196__I _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4709__I _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7169_ _1081_ _1070_ _1634_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7787__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7787__B2 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6924__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4444__I _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A1 _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6762__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4773__A1 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5275__I _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7490__I _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6278__A1 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4619__I _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5878__C _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _0469_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6202__A1 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6753__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6540_ _1807_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6471_ _1933_ _1934_ _1931_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6505__A2 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7702__A1 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ net35 _3557_ _3472_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5422_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8141_ _2827_ _3442_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5353_ _0882_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4304_ _3875_ _3884_ _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8072_ _0395_ _0422_ _3423_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_102_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4819__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7023_ _1390_ _1416_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4529__I _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5492__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__A1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8430__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5244__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _3256_ _3284_ _3291_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4264__I _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7856_ _1131_ _1594_ _3247_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8194__A1 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6807_ _4049_ _2114_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7787_ _1473_ _1423_ _1389_ _3189_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6744__A2 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _0595_ _0593_ _0597_ _0349_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7941__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _2167_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _0308_ _2120_ _2129_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8408_ _0685_ _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8339_ _3081_ _3680_ _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8249__A2 _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6919__I _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5180__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7457__B1 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4439__I _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6680__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5979__B _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8074__C _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__A1 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6735__A2 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6603__B _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4746__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8488__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_17_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6499__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6829__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5171__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7999__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8660__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8412__A2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5226__A2 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6423__A1 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _1488_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6974__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7710_ _4157_ _2037_ _2544_ _3116_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4922_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8690_ _0167_ clknet_leaf_0_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8176__A1 _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7641_ _2893_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4853_ _0433_ _0427_ _0450_ _0453_ _0426_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7395__I as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__B _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7923__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4812__I _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7572_ _2662_ _2970_ _2972_ _2885_ _2983_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7328__C _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4784_ _0383_ _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6454_ _1916_ _1936_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5405_ _0924_ as2650.stack\[3\]\[14\] as2650.stack\[2\]\[14\] _0941_ _0995_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _0390_ _1759_ _1868_ _1658_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8124_ net32 _3445_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7439__B1 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5336_ as2650.r123\[0\]\[1\] _0860_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8100__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8055_ _3316_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5267_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6662__A1 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7006_ _1357_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5465__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ _0770_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8403__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6414__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5217__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5768__A3 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7908_ as2650.stack\[3\]\[13\] _1249_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7839_ as2650.stack\[6\]\[0\] _1602_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4728__A1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__B2 _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5039__B _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7142__A2 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8683__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4900__A1 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6653__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5456__A2 _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7905__A1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A1 _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5392__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5392__B2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7133__A2 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8330__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8330__B2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A1 _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__I _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6170_ _4137_ _1652_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5121_ _4226_ _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5447__A2 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6644__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5052_ _0650_ _0578_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7611__C _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6508__B _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8397__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6947__A2 _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4958__A1 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8742_ _0219_ clknet_leaf_39_wb_clk_i as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5954_ _4092_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8149__A1 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__C _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4905_ _0431_ _0438_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8673_ _0150_ clknet_leaf_17_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5885_ _3954_ _1398_ _1402_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8556__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7624_ _2639_ _3033_ _2694_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4836_ _0353_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7372__A2 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7555_ as2650.pc\[9\] _1157_ _2902_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5383__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6506_ as2650.r123_2\[2\]\[6\] _1910_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7486_ _2523_ _2898_ _2900_ _2633_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8321__A1 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4698_ _4105_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7074__B _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6437_ _1918_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6883__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6368_ _1850_ _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8107_ _0543_ _0518_ _3457_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5319_ _0861_ _0914_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6299_ _1745_ _1784_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6635__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ _3326_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8388__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6938__A2 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7363__A2 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7763__I _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5913__A3 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8312__A1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5126__A1 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6874__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6874__B2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8076__B1 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5429__A2 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4627__I _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7003__I _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8379__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__A3 _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5458__I _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_32_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5670_ _1220_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5365__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ _4200_ _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7673__I _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7340_ _2531_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7606__C _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4552_ _3994_ _4132_ _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8303__A1 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7106__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8303__B2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7271_ _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4483_ _4063_ _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5668__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _4140_ _1708_ _3937_ _1691_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6153_ _1645_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4340__A2 _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6617__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5104_ _0494_ _0383_ _0537_ _0676_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_98_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6084_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6093__A2 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6632__A4 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6986_ _2356_ _1327_ _2415_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8725_ _0202_ clknet_leaf_74_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5937_ _0603_ _1376_ _1325_ _1384_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4272__I _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8656_ _0133_ clknet_leaf_71_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _3867_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7345__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7607_ _3017_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5356__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4819_ _4044_ _0386_ _0387_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8587_ _0064_ clknet_leaf_32_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6699__A4 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5799_ _1288_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7538_ _2662_ _2950_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6420__C _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7469_ _2614_ _2880_ _2883_ _2264_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput13 net50 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5659__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput35 net35 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_66_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7281__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8721__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5987__B _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A2 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7584__A2 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4398__A2 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5278__I _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6544__B1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6330__C _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8064__A3 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7272__A1 _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8273__B _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7024__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6840_ _2280_ _2282_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6771_ _1046_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8510_ _1297_ _0462_ _3816_ _3832_ _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5722_ _1232_ _1250_ _1255_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7327__A2 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8441_ _1058_ _3138_ _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5653_ _1137_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5916__I _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5889__A2 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _3981_ _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8372_ _3699_ _3707_ _3708_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5584_ _1013_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7323_ _1100_ _2699_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4535_ _4055_ _4061_ _4114_ _4115_ _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4561__A2 _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6838__A1 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7254_ _2667_ _2670_ _2672_ _2673_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_4466_ _4046_ _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6205_ _4050_ _1691_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4313__A2 as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8744__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5510__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ _2600_ _2602_ _2605_ _1614_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6853__A4 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _3968_ _3974_ _3977_ _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _1634_ _1629_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4864__A3 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4267__I _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ _1089_ _1576_ _1581_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5018_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6415__C _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _2375_ _2235_ _2399_ _2346_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_74_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8708_ _0185_ clknet_leaf_36_wb_clk_i as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8515__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8639_ _0116_ clknet_leaf_66_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__A2 _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8358__B _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6657__I _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4304__A2 _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5501__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6606__B _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7557__A2 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8617__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8506__A1 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6780__A3 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7437__B _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8767__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6995__C _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4320_ _3888_ _3899_ _3900_ _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7493__A1 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6296__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6567__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5471__I _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4697__I3 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7245__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__B1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7796__A2 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7941_ _1234_ _3298_ _3301_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6516__B _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7872_ as2650.stack\[5\]\[12\] _3252_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7548__A2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _1503_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6754_ _2199_ _1857_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8450__C _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5705_ as2650.stack\[2\]\[5\] _1235_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6685_ as2650.addr_buff\[7\] _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4782__A2 _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7066__C _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5636_ _1163_ _1200_ _1201_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8424_ _0605_ _0611_ _3739_ _1976_ _3754_ _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7720__A2 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8355_ net43 _3688_ _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5567_ _1103_ _1136_ _1143_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7861__I _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7306_ _2635_ _2685_ _2724_ _2630_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4518_ _4098_ _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8286_ _3330_ _3630_ _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8178__B _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5498_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7237_ _1512_ _4085_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6287__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7484__A1 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4449_ _4020_ _4008_ _4022_ _4026_ _4029_ _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_132_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7168_ _1069_ _2292_ _1081_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7236__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6119_ _1606_ _1613_ _1619_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7099_ _2520_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7787__A2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7101__I _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4470__A1 _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A2 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6940__I _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5556__I _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6278__A2 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6202__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7950__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4370__I _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _1915_ _1937_ _1951_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5421_ _3956_ _1007_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5713__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8140_ _2461_ _3489_ _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5352_ _0924_ as2650.stack\[3\]\[10\] as2650.stack\[2\]\[10\] _0920_ _0946_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_126_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4303_ _3883_ _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8071_ _3394_ _3421_ _3422_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5283_ _0876_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_82_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7022_ _1366_ _2450_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4819__A3 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7218__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7769__A2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5324__S0 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6441__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7924_ as2650.stack\[7\]\[11\] _3288_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7855_ as2650.stack\[6\]\[7\] _1591_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8194__A2 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6806_ _4048_ _1314_ _2089_ _2113_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_4998_ _0586_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7786_ _1509_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7941__A2 _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6737_ net23 _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4280__I _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6668_ _2128_ _2126_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8407_ _1428_ _3737_ _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5619_ _1186_ _1073_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7805__B _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6599_ as2650.r123_2\[0\]\[6\] _2045_ _2030_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8338_ _3675_ _2228_ _3679_ _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__A2 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8249__A3 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7457__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8269_ net37 _3557_ _3614_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6504__I0 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7457__B2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6000__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6680__A2 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6432__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6670__I _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7932__A2 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5943__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__I _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6499__A2 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7160__A3 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5171__A2 _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_57_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7006__I _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7999__A2 _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6845__I _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8265__C _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6959__B1 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6423__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5970_ _1487_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _3858_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4985__A2 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8176__A2 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8712__D _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4852_ _0357_ _0452_ _0358_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7640_ _3024_ _3049_ _2992_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6187__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7923__A2 _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7571_ _2834_ _2978_ _2982_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4783_ _0311_ _0328_ _0381_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5934__A1 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _3849_ _1711_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7687__A1 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6453_ _1931_ _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5404_ _0920_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6384_ _1860_ _1866_ _1867_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8123_ _3408_ _3471_ _3473_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7439__A1 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7439__B2 _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5335_ _0859_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8100__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8054_ _3343_ _3405_ _3406_ _3224_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5266_ _3914_ _0850_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7005_ _2164_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6662__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5197_ _0773_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8175__C _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4275__I _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__A2 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__A1 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__A4 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _3258_ _1252_ _3279_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8167__A2 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6178__A1 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7838_ _2068_ _3130_ _3237_ _3224_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_93_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__A2 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7769_ _1530_ _4223_ _3172_ _3120_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7678__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7535__B _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6653__A2 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7850__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4664__A1 _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4416__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8158__A2 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7905__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7381__A3 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5392__A2 as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7669__A1 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8330__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _0682_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6644__A2 _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5051_ _0478_ _0480_ _0577_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8397__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4407__A1 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8741_ _0218_ clknet_leaf_35_wb_clk_i as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5953_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _0427_ _0452_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8672_ _0149_ clknet_leaf_17_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5884_ _1400_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7623_ as2650.pc\[12\] _3032_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5907__A1 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4835_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4766_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5383__A2 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6580__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7554_ _2965_ _2772_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6505_ _1808_ _1985_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7485_ _2867_ _2899_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4697_ as2650.r123\[1\]\[3\] as2650.r123\[0\]\[3\] as2650.r123_2\[1\]\[3\] as2650.r123_2\[0\]\[3\]
+ _3857_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8030__I _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ _1884_ _1885_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6332__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6883__A2 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6367_ _1779_ _1802_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8085__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5318_ _4153_ _0867_ _0869_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8106_ _3455_ _3456_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7802__C _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6298_ _1748_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6635__A2 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7832__A1 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5249_ as2650.r123\[1\]\[7\] _4253_ _0845_ _4149_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8037_ _1518_ _3383_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4646__A1 _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8388__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4934__S _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6399__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4949__A2 _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5829__I _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7348__B1 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8650__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6571__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8312__A2 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8076__A1 _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8076__B2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8379__A2 _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5062__A1 _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4643__I _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _3865_ _4141_ _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_72_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4551_ _3943_ _4019_ _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5474__I _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8303__A2 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7270_ as2650.pc\[2\] net7 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4482_ net5 _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5117__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _1707_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8067__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6152_ as2650.r123\[3\]\[2\] _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4340__A3 as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5103_ _0588_ _0619_ _0633_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6617__A2 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7814__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A1 _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _0628_ _0630_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8523__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6985_ _2410_ _2412_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8025__I _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8724_ _0201_ clknet_leaf_77_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5936_ _4229_ _1428_ _1431_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__8673__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4800__A1 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8655_ _0132_ clknet_leaf_71_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5867_ _1384_ _1319_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7606_ _2781_ _2996_ _3008_ _2732_ _2592_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5356__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _0417_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_8586_ _0063_ clknet_leaf_32_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5798_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7537_ _2125_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4749_ _4020_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6305__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7468_ _2396_ _2881_ _2094_ _2142_ _2882_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_68_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput14 net14 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput25 net25 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6419_ _1899_ _1901_ _1684_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput36 net36 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7399_ _2624_ as2650.stack\[5\]\[6\] as2650.stack\[4\]\[6\] _2625_ _2815_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7805__A1 _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6943__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5831__A3 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8230__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6792__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A3 _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8297__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A2 _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7723__B _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8049__A1 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7014__I _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8696__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7024__A2 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5469__I _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4373__I _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6783__A1 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6770_ _1044_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7980__B1 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5721_ as2650.stack\[3\]\[1\] _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8720__D _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8440_ _2146_ _0444_ _1368_ _0863_ _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6535__A1 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _1078_ _1200_ _1210_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4603_ _3995_ _4028_ _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8371_ net19 _3704_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5889__A3 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5583_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8288__A1 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7322_ _2732_ _2737_ _2739_ _2565_ _2392_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4534_ _4038_ _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6838__A2 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7253_ _2534_ as2650.stack\[3\]\[2\] as2650.stack\[2\]\[2\] _2535_ _1021_ _2673_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4465_ _4032_ _4045_ _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5932__I _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4849__A1 _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6204_ _1673_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7184_ _1516_ _2604_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7352__C _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4313__A3 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4396_ _3975_ _3976_ _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4548__I _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6135_ _1633_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ as2650.stack\[5\]\[1\] _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8460__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4283__I _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6774__A1 _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6968_ _2380_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5577__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8707_ _0184_ clknet_leaf_37_wb_clk_i as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5919_ _4008_ _4027_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6899_ _2335_ _0444_ _1455_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8515__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8630__D _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8638_ _0115_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8569_ _0046_ clknet_leaf_46_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8279__A1 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4458__I _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8451__A1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8203__A1 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5289__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6765__A1 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6517__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7190__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5752__I _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8442__B2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__A1 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7940_ as2650.stack\[7\]\[2\] _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7871_ _1188_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5008__A1 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5008__B2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6822_ net26 _1349_ _2265_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6756__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5559__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6753_ _4252_ _2194_ _2201_ _2203_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5704_ _1119_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6684_ _1506_ _2123_ _2140_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4782__A3 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5148__B _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8423_ _3741_ _3742_ _3753_ _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5635_ as2650.stack\[2\]\[14\] _1195_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8711__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8354_ _3684_ _4223_ _3693_ _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5566_ as2650.stack\[1\]\[3\] _1140_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5731__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8459__B _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7305_ _0880_ _2720_ _2723_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4517_ as2650.r0\[7\] _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8285_ _3628_ _3629_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5497_ _3986_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8178__C _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7236_ net7 _4216_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4448_ _4021_ _4027_ _4028_ _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4379_ _3959_ _3892_ _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7167_ _2548_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6118_ _1609_ _1617_ _1618_ _4139_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7236__A2 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ _2519_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ _1563_ _1334_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6995__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A2 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8213__I _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5722__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8424__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8424__B2 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7720__C _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6986__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8734__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5410__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7163__A1 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7962__I _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _3973_ _0530_ _0862_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_51_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5351_ _0942_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4302_ _3879_ _3882_ _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5282_ as2650.psu\[2\] _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8070_ _0306_ _0325_ _0330_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_142_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ _3893_ _1028_ _2302_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5229__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6977__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5324__S1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7923_ _3254_ _3284_ _3290_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__A2 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6729__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7854_ _1127_ _1594_ _3246_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6805_ _1610_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7785_ _3123_ _1474_ _1408_ _2176_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4997_ _0447_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6736_ _2174_ _2178_ _2188_ _1338_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6667_ as2650.addr_buff\[2\] _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8406_ as2650.holding_reg\[7\] _0595_ _3736_ _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5618_ _0568_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6901__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6901__B2 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ _2061_ _2063_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8337_ _2092_ _3094_ _3677_ _3678_ _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5549_ _1129_ _1004_ _1110_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8268_ _2166_ _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5468__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7219_ _2564_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8199_ net34 net33 _3474_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8607__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8406__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4443__A2 _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7393__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7715__C _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5459__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26_wb_clk_i clknet_opt_2_1_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6959__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6959__B2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7620__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6861__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _3971_ _0382_ _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7384__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6187__A2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7570_ _2611_ _2968_ _2981_ _2654_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4782_ _4032_ _4091_ _4221_ _0301_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _1859_ _1990_ _1999_ _1713_ _2000_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_53_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7136__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7692__I _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7687__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6452_ _1933_ _1934_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5403_ _0921_ as2650.stack\[1\]\[14\] as2650.stack\[0\]\[14\] _0943_ _0993_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6383_ _0422_ _1687_ _1697_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8122_ net32 _3317_ _3472_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5334_ _4198_ _0917_ _0868_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8053_ net30 _3342_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5265_ _0859_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _2408_ _2432_ _2433_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5196_ _0780_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5870__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__A2 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6771__I _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7906_ as2650.stack\[3\]\[12\] _3275_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7837_ _3227_ _3236_ _3101_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5387__I as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7375__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4291__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7768_ _3116_ _2724_ _3170_ _2038_ _3171_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6719_ _2170_ _2171_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7699_ _2850_ _3104_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7678__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5689__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7107__I _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7551__B _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6946__I _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5850__I _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6102__A2 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7850__A2 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4664__A2 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4466__I _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7602__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4416__A2 _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7366__A1 _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5297__I _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7669__A2 _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7017__I _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6856__I _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5050_ _3993_ _0611_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_61_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5852__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4655__A2 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4407__A2 _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__A1 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8723__D _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8740_ _0217_ clknet_leaf_49_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5952_ _1385_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4903_ _0495_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8671_ _0148_ clknet_leaf_21_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5883_ _3847_ _1399_ _1350_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_90_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7357__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7622_ _2993_ _2994_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4834_ _3971_ _0310_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5907__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7553_ as2650.pc\[10\] _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4765_ _0366_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _1976_ _1984_ _1695_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7484_ _2573_ _2896_ _2696_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4696_ _3853_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8321__A3 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _1840_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4343__A1 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6366_ _1781_ _1801_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8467__B _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8105_ _0394_ _0421_ _3394_ _3421_ _3422_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _0871_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8085__A2 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6297_ _0783_ _1782_ _1741_ _1739_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_88_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8036_ _3386_ _3387_ _3388_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5248_ _0820_ _0823_ _0844_ _4162_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7832__A2 _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4646__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4286__I _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5179_ _0661_ _0774_ _0775_ _0748_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_112_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8388__A3 _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7596__A1 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6715__B _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7348__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6020__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5845__I _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7520__A1 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7520__B2 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8076__A2 _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4637__A2 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5834__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__A1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4550_ _3957_ _4130_ _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _4059_ _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5117__A3 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4325__A1 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6220_ _3931_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8287__B _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8067__A2 _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _1644_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_41_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5102_ _0676_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _1133_ _1151_ _1573_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7814__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A2 _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _4105_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7578__A1 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6984_ _2344_ _2413_ _2398_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6250__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8723_ _0200_ clknet_leaf_77_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5935_ _4176_ _1433_ _1436_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_80_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8654_ _0131_ clknet_leaf_71_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5866_ _4012_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_90_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7605_ _1532_ _3011_ _3015_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _4242_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8585_ _0062_ clknet_leaf_34_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5797_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6553__A2 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7536_ _2552_ _2920_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4564__A1 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _4163_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7467_ _2612_ _2867_ _1605_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4679_ _4257_ _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4316__A1 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6418_ _1900_ _1683_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput15 net15 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput26 net26 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7398_ _2812_ _2813_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput37 net37 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8628__D _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6349_ _1788_ _1833_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6069__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8019_ _2316_ _3368_ _3372_ _2299_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7569__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8216__I _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8230__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6792__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7276__B _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7741__A1 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4555__A1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__I _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5807__A1 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6783__A2 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7980__A1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ _1251_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ as2650.stack\[0\]\[14\] _1066_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5485__I _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6535__A2 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__A1 _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _4175_ _4181_ _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8370_ _3700_ _1474_ _3706_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5582_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7321_ _1108_ _2738_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4533_ _4062_ _4113_ _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8288__A2 _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7252_ _0893_ _2671_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6838__A3 _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ _4042_ _4044_ _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6203_ _1689_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7183_ _2603_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4395_ as2650.idx_ctrl\[0\] _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_98_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6134_ _1052_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6065_ _1577_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8460__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5016_ net1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8640__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__A1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _2396_ _4204_ _2397_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6774__A2 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7971__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5918_ _0428_ _0430_ _1435_ _0343_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8706_ _0183_ clknet_leaf_37_wb_clk_i as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6898_ _2289_ _2253_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8515__A3 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8637_ _0114_ clknet_leaf_61_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5849_ _1364_ _1320_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5395__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6526__A2 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7723__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4537__A1 _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8568_ _0045_ clknet_leaf_45_wb_clk_i as2650.stack\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7519_ _2852_ _2921_ _2932_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8499_ _2357_ _3819_ _4097_ _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6954__I _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8451__A2 _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6462__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4474__I _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8203__A2 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8390__B _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6765__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7718__C _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6517__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7190__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8663__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7245__A3 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7870_ _3256_ _3249_ _3257_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6205__A1 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _2264_ _2149_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7953__A1 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7695__I _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6752_ as2650.r123\[2\]\[1\] _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ _1239_ _1240_ _1241_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _2139_ _2119_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7705__A1 _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4782__A4 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6104__I _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8422_ _3743_ _3751_ _3752_ _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5634_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8353_ _1094_ _3685_ _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5565_ _1097_ _1136_ _1142_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7304_ _0893_ _2721_ _2722_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4516_ as2650.psl\[3\] _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8284_ net37 net51 _3567_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8130__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5496_ _3884_ _1008_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7235_ _2651_ _2653_ _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4447_ _3870_ _4012_ _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7166_ _1617_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4378_ as2650.cycle\[3\] _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6117_ _1562_ _1332_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _2259_ _2506_ _2510_ _2518_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_115_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6048_ _1561_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4294__I _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8197__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7944__A1 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7999_ _1556_ _3351_ _3352_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6949__I _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8686__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4930__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__A1 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8424__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A1 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6986__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8188__A1 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7935__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4932__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5410__A2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__I0 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6859__I _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _0921_ as2650.stack\[1\]\[10\] as2650.stack\[0\]\[10\] _0943_ _0944_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_138_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8112__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4301_ _3880_ _3881_ _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5281_ _0872_ _0873_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _2441_ _2445_ _2447_ _2448_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5477__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8726__D _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6426__A1 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5229__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4988__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7922_ as2650.stack\[7\]\[10\] _3288_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7853_ as2650.stack\[6\]\[6\] _1591_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8559__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6729__A2 _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5938__I _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6804_ _2104_ _2247_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__I _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7784_ _3153_ _3186_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4996_ _0447_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6735_ _1323_ _2182_ _2185_ _2187_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6666_ _4225_ _2120_ _2127_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8351__A1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8405_ _0595_ _1456_ _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5617_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6597_ _0967_ _2062_ _2048_ _0986_ _2054_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6901__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8336_ _1463_ _1450_ _2182_ _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5548_ as2650.pc\[7\] _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8267_ _3607_ _3612_ _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5479_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5468__A2 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6665__A1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7218_ _1092_ _2637_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8198_ _3537_ _3538_ _3544_ _3545_ _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8406__A2 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7149_ _2524_ _2527_ _2529_ _2545_ _2570_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7090__A1 _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7393__A2 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout50 net13 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6679__I _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5459__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6959__A2 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7081__A1 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8701__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_66_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7908__A1 as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _0429_ _3971_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7384__A2 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6187__A3 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6041__C1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _0381_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6520_ as2650.r123_2\[2\]\[7\] _1910_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8333__A1 _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7136__A2 _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _1834_ _1889_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__I as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ as2650.stack\[7\]\[14\] as2650.stack\[4\]\[14\] as2650.stack\[5\]\[14\] as2650.stack\[6\]\[14\]
+ _0938_ _0939_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6382_ _0391_ _1663_ _1864_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8121_ _2166_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5333_ _0871_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6647__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8052_ _1093_ _3377_ _3404_ _2331_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7003_ _2276_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5195_ _0781_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7072__A1 _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5622__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7905_ _3256_ _3273_ _3278_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4572__I _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7836_ _1457_ _3137_ _3228_ _3235_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4979_ _0467_ _0481_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7767_ _0472_ _3156_ _4207_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6718_ _1031_ _3879_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8324__A1 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7698_ _2402_ _4047_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _2110_ _2111_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7678__A3 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6886__A1 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5689__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8319_ net39 _3645_ _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4747__I _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8219__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8724__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7123__I _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7063__A1 as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6810__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4482__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6023__C1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7366__A2 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5377__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4424__I0 _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__B2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8315__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5129__A1 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5246__C _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6629__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__I _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5852__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7968__I _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7054__A1 _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5604__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6801__A1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7189__B _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ _1411_ _1468_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5488__I _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4392__I _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _0358_ _0489_ _0501_ _0349_ _4170_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8670_ _0147_ clknet_leaf_7_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5882_ _1048_ _1399_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7357__A2 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7621_ _2567_ _3030_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5368__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4833_ as2650.holding_reg\[2\] _3970_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5907__A3 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7552_ _2809_ _2963_ _2964_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4764_ as2650.r123\[0\]\[2\] as2650.r123_2\[0\]\[2\] _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6503_ _0706_ _1809_ _1983_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7483_ _2527_ _2867_ _2874_ _2875_ _2897_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4695_ _4101_ _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6868__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6434_ _0612_ _1837_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6365_ _1848_ _1849_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5540__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8747__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__A2 _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8467__C _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8104_ _0394_ _0421_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5316_ _0882_ _0888_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _0532_ _0568_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7293__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8035_ _3386_ _3387_ _3349_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5247_ _0831_ _0843_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5178_ _0293_ _0471_ _0567_ _4214_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8483__B _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6782__I _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7348__A2 _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7819_ _1485_ _1507_ _3219_ _2592_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8799_ _0276_ clknet_leaf_34_wb_clk_i as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6020__A2 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7546__C _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7118__I _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6022__I _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7520__A2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5861__I _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7284__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6087__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__A2 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6692__I _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__B _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__A2 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__B1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4940__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6011__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4480_ _4060_ _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4325__A2 _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ as2650.r123\[3\]\[1\] _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5101_ _0536_ _0620_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4387__I _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _1131_ _1584_ _1589_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ as2650.r123\[1\]\[6\] as2650.r123\[0\]\[6\] as2650.r123_2\[1\]\[6\] as2650.r123_2\[0\]\[6\]
+ _3845_ _3855_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6816__B _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7027__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_10_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5589__A1 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6983_ _1040_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8722_ _0199_ clknet_leaf_77_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ _1448_ _1449_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5865_ _1364_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8653_ _0130_ clknet_leaf_75_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5946__I _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7604_ _2379_ _2995_ _3014_ _2422_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4816_ _4043_ _3935_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5796_ _1313_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8584_ _0061_ clknet_leaf_34_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5761__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _4013_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7535_ _2905_ _2947_ _2858_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4564__A2 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7466_ _2384_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4678_ _4197_ _4053_ _4157_ _4257_ _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_135_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6417_ _0398_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7382__B _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5513__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7397_ _1115_ _2773_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput16 net16 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput27 net27 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput38 net38 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6348_ _4098_ _0568_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6279_ _1556_ _1670_ _1764_ _1667_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8018_ _1082_ _3337_ _3371_ _2304_ _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7018__A1 _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6017__I _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8518__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7276__C _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7741__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7257__A1 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5807__A2 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5363__S0 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7009__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8206__B1 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__A1 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8509__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7980__A2 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7467__B _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8592__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__I _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _1078_ _1194_ _1209_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _4033_ _4027_ _4011_ _4017_ _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__A2 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _1011_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5743__A1 as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7320_ _1100_ _2684_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ _4075_ _4096_ _4111_ _4112_ _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8298__B _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7251_ _0899_ as2650.stack\[1\]\[2\] as2650.stack\[0\]\[2\] _0895_ _2671_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4463_ _4043_ _3935_ _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6202_ _4141_ _1673_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7182_ _1036_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ as2650.idx_ctrl\[1\] _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_98_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _1629_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__A2 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _1076_ _1576_ _1579_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _0499_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4845__I _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7420__A1 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6966_ _2078_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7971__A2 _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8705_ _0182_ clknet_leaf_37_wb_clk_i as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5917_ _1434_ _4175_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4785__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6897_ _2071_ _2335_ _2336_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_107_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4580__I _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8636_ _0113_ clknet_3_5_0_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8515__A4 _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5848_ _1365_ _1342_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6526__A3 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4537__A2 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5734__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8567_ _0044_ clknet_leaf_46_wb_clk_i as2650.stack\[0\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5779_ as2650.psl\[6\] _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7518_ _2588_ _2925_ _2930_ _2931_ _2854_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7824__C _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8498_ _3820_ _3823_ _2992_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7449_ _2863_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6462__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4755__I _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6970__I _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__A2 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4665__I _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7650__A1 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A1 _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6205__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7402__A1 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6820_ _2263_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7402__B2 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _2196_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ as2650.stack\[2\]\[4\] _1235_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6682_ _3935_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8421_ _0489_ _0509_ _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4519__A2 _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ as2650.pc\[14\] _1179_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8352_ _3682_ _3691_ _3692_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5564_ as2650.stack\[1\]\[2\] _1140_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7469__A1 _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4515_ _4078_ _4092_ _4095_ _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7303_ _2534_ as2650.stack\[3\]\[3\] as2650.stack\[2\]\[3\] _2540_ _2536_ _2722_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_8283_ net38 _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5495_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7216__I _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6120__I _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7234_ _1296_ _2546_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4446_ _4010_ _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6141__A1 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7165_ _2215_ _2247_ _2585_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4377_ _3896_ _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6116_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7096_ _1363_ _2511_ _2517_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4575__I _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6047_ _1538_ _1563_ _1324_ _1351_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4455__A1 _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8491__B _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7819__C _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ _4063_ _4123_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7944__A2 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4758__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _2308_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8619_ _0096_ clknet_leaf_52_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7835__B _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6380__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4930__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6132__A1 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7570__B _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6965__I _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__A2 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5090__B _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7632__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8188__A2 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6199__A1 _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7729__C _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7935__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7699__A1 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5549__I1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8360__A2 _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8630__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7036__I _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4300_ as2650.cycle\[0\] _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6123__A1 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5280_ _0872_ _0874_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8780__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4685__B2 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6426__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7623__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4395__I as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4437__A1 _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7921_ _3251_ _3284_ _3289_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4988__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7852_ _1120_ _1594_ _3245_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6803_ _2241_ _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5937__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7783_ _1531_ _1900_ _3185_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4995_ as2650.holding_reg\[5\] _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6115__I _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6734_ _2183_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7655__B _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6665_ _2125_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5954__I _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8404_ _3717_ _3728_ _3735_ _2435_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5616_ as2650.pc\[12\] _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6596_ _0985_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8335_ _4139_ _3964_ _2237_ _3676_ _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5547_ _1105_ _1127_ _1128_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8266_ _1166_ _3377_ _3608_ _3611_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5478_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8486__B _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6665__A2 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4429_ _4009_ _4006_ _3980_ _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7217_ _1080_ _1068_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8197_ _2396_ _3454_ _2485_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7148_ _1636_ _2563_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7614__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7079_ net4 _1401_ _2498_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7090__A2 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7917__A2 _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout51 net36 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8653__CLK clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__I _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6353__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__A2 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8396__B _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4667__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7081__A2 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4943__I _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7908__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5919__A1 _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__B1 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6041__C2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6187__A4 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4780_ _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6592__A1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7475__B _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8333__A2 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6450_ _1878_ _1932_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5401_ _0727_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6381_ _0392_ _1683_ _1684_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8120_ _2730_ _3377_ _3470_ _2331_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5332_ _0918_ _0919_ _0923_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8097__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8051_ _3168_ _3400_ _3403_ _3126_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6647__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _4128_ _0857_ _0858_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_130_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4658__A1 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7002_ _2319_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5194_ _0745_ _0784_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_99_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__CLK clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5014__I _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5083__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5949__I _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7904_ as2650.stack\[3\]\[11\] _3275_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7369__C _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8676__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8021__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8021__B2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7835_ _1641_ _2176_ _2177_ _3234_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6032__B1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6583__A1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7766_ _1554_ _4016_ _3110_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4978_ _0467_ _0481_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6717_ _1335_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4802__B _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7697_ _3103_ _4124_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8324__A2 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6648_ _3928_ _3890_ _3929_ _2073_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6335__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6886__A2 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6579_ _0871_ _1653_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4897__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8318_ _3591_ _3660_ _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7835__A1 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8249_ _2121_ _3576_ _3578_ _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4649__A1 as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7063__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5859__I _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__B1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__C2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4424__I1 _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7295__B _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8315__A2 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5129__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6326__A1 _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8079__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7742__C _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6629__A2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4938__I _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7826__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7314__I _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8699__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A2 _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5065__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6801__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5950_ _1467_ _0813_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _0447_ _0499_ _0500_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ _3947_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7620_ _3028_ _3029_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_94_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _4170_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7551_ _2952_ _2633_ _2938_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4763_ as2650.psl\[4\] _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _0709_ _1810_ _1697_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7482_ _2884_ _2895_ _2896_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4694_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _3854_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6868__A2 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6433_ _1890_ _1893_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6364_ _1824_ _1825_ _1847_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5540__A2 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8103_ _3083_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7817__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5315_ _0894_ _0902_ _0909_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6295_ _1735_ _1751_ _1780_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8490__A1 _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8034_ _0304_ _0337_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7293__A2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5246_ _0839_ _0841_ _0842_ _0609_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5177_ as2650.r0\[3\] _0566_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8242__A1 _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8242__B2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4583__I _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8055__I _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6504__S _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7818_ _3143_ _4110_ _3218_ _1470_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7827__C _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8798_ _0275_ clknet_leaf_35_wb_clk_i as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7749_ as2650.overflow _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7808__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7284__A2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8481__A1 _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5295__A1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4694__S _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8393__C _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6795__A1 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5100_ _0609_ _0678_ _0697_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_98_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ as2650.stack\[5\]\[7\] _1586_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8472__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _4102_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7027__A2 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__I _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5038__A1 _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6786__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6982_ _2403_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5589__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7983__B1 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8721_ _0198_ clknet_leaf_77_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _1450_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_50_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8652_ _0129_ clknet_leaf_72_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6538__A1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7735__B1 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7603_ _2547_ _3013_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4815_ _0391_ _4062_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8583_ _0060_ clknet_leaf_59_wb_clk_i as2650.r123_2\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5795_ _3879_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7219__I _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8714__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7534_ _2906_ _2941_ _2946_ _2915_ _2916_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_72_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4746_ _0343_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5761__A2 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4564__A3 _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7663__B _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7465_ _2876_ _2879_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4677_ _4256_ _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6416_ _0540_ _1668_ _1898_ _1680_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5513__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7396_ _2811_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput17 net17 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput28 net28 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput39 net39 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6347_ _4098_ _0472_ _1186_ _0626_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8463__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _1763_ _1669_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8494__B _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8017_ _2418_ _2598_ _3332_ _3370_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5229_ _0824_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7018__A2 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5029__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__B1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8518__A2 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6461__C _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A1 _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7129__I _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6968__I _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6701__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5504__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4488__I _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7257__A2 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5268__A1 _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__B1 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5821__B _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5363__S1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7009__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8206__A1 _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8206__B2 _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__A2 _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6208__I _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6768__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5112__I _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5440__A1 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8737__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8509__A2 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _3995_ _4020_ _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5580_ _1151_ _1063_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5743__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6878__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _4094_ _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7496__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7250_ as2650.stack\[6\]\[2\] _2668_ _1015_ _2669_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4462_ as2650.addr_buff\[5\] _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6201_ _4054_ _1663_ _1681_ _1685_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7181_ _2558_ _2601_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4393_ _3973_ _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8445__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _1626_ _1627_ _1631_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ as2650.stack\[5\]\[0\] _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7502__I _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6759__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7420__A2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6223__A3 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _1562_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8704_ _0181_ clknet_leaf_17_wb_clk_i as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _4130_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6281__C _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4785__A3 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__A2 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6896_ _4054_ _2146_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8635_ _0112_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5847_ _3875_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7184__A1 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8566_ _0043_ clknet_leaf_45_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5734__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5778_ _0529_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7393__B _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7517_ _2654_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4729_ _0325_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8497_ _3822_ _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7448_ as2650.pc\[7\] _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7379_ _2442_ _2774_ _2779_ _4144_ _2795_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8436__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__A1 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7411__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5973__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7175__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__A2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8399__B _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8427__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7650__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A2 _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _2199_ _1804_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ _1229_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6681_ _2136_ _2123_ _2138_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8420_ _0452_ _0455_ _3744_ _3749_ _3750_ _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5632_ _1197_ _1073_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6913__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8351_ net42 _3688_ _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5563_ _1089_ _1136_ _1141_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7302_ _0899_ as2650.stack\[1\]\[3\] as2650.stack\[0\]\[3\] _0895_ _2721_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7469__A2 _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4514_ _4094_ _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8282_ _3410_ _3626_ _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5494_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7233_ _2300_ _2646_ _2652_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4445_ _4025_ _4011_ _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7164_ _2355_ _2584_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4376_ _3952_ _3956_ _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5461__B _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ _1615_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8328__I _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ _2091_ _2230_ _2516_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _1562_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5652__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5404__A1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ _4006_ _4166_ _4248_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5687__I _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6948_ _1392_ _2247_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6879_ _2319_ _3904_ _2079_ _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8618_ _0095_ clknet_leaf_56_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7835__C _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8549_ _0026_ clknet_leaf_52_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7570__C _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5891__A1 _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8582__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4766__I _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7632__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6930__B _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7148__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6221__I _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4382__A1 _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6123__A2 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7320__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7480__C _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5882__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4685__A2 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__I _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7920_ as2650.stack\[7\]\[9\] _3288_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6824__C _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7851_ as2650.stack\[6\]\[5\] _3241_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7387__A1 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6802_ _2242_ _0810_ _2245_ _1302_ _4132_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5300__I _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7782_ _1186_ _2286_ _3184_ _1495_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4994_ _0588_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5937__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6733_ _3903_ _1289_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _2118_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8403_ _3671_ _0511_ _3728_ _3734_ _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5615_ _1155_ _1182_ _1183_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6595_ _1948_ _2028_ _2034_ _2060_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8334_ _4056_ _2155_ _1389_ _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5546_ as2650.stack\[0\]\[6\] _1121_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8265_ _2952_ _3495_ _3497_ _3610_ _2522_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6114__A2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5970__I _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ _1011_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7311__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8486__C _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7216_ _2635_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4428_ as2650.holding_reg\[0\] _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8196_ _3541_ _3542_ _3543_ _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5873__A1 _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8058__I _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7147_ _2524_ _2565_ _2568_ _2426_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4359_ _3872_ _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7614__A2 _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7078_ _2068_ _2498_ _2500_ _1401_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5625__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6029_ net3 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7378__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4535__B _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5210__I _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6050__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__B2 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net33 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7550__A1 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7550__B2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4364__A1 _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7581__B _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__B2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7853__A2 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4667__A2 as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7369__A1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7369__B2 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_90 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_127_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__B2 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7756__B _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7541__A1 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5147__A3 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4355__A1 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ as2650.r123\[0\]\[6\] _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6380_ _0614_ _1668_ _1863_ _1680_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_75_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5331_ _0918_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8097__A2 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8050_ _1093_ _3337_ _3402_ _2304_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5262_ _0848_ _4148_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7001_ _2159_ _2416_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5855__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _0785_ _0786_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_64_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5607__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6280__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7903_ _3254_ _3273_ _3277_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__A2 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8021__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7834_ _1497_ _3233_ _1469_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6032__A1 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6032__B2 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7765_ _3164_ _0456_ _3165_ _3166_ _3168_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4977_ _0574_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6583__A2 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7780__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8341__I _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6716_ _3870_ _2165_ _2169_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7385__C _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7696_ _2322_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6647_ _2108_ _2109_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7532__A1 _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6335__A2 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _1821_ _2027_ _2030_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8317_ _2134_ _3641_ _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8088__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ as2650.stack\[0\]\[4\] _1090_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8248_ net37 _3593_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7835__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4649__A2 _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8179_ _3509_ _3527_ _2333_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7599__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7063__A3 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6271__A1 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8620__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6023__B2 _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8770__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7771__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4424__I2 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7295__C _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4337__A1 _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8079__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__A2 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5837__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A3 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8251__A2 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5065__A2 _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6801__A3 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ _0485_ _4184_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _1044_ _1294_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7762__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7550_ _2941_ _2948_ _2962_ _2935_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4762_ _0333_ _0338_ _0363_ _4162_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_92_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ _1977_ _1981_ _1686_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7481_ _2732_ _2880_ _2867_ _2781_ _2592_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__7514__A1 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ _0294_ _3859_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6432_ _1853_ _1856_ _1913_ _1914_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6363_ _1824_ _1825_ _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8110__B _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8102_ _3383_ _3451_ _3452_ _3348_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5314_ _0881_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7817__A2 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6294_ _1738_ _1750_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8033_ _3352_ _3384_ _3385_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_130_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5245_ as2650.holding_reg\[7\] _0433_ _4110_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8490__A2 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8643__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ _0771_ _0756_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6565__B _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8242__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6253__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5056__A2 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6284__C _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8793__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6005__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7202__B1 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7817_ _1477_ _0540_ _3217_ _1467_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_40_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4813__B _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8797_ _0274_ clknet_leaf_38_wb_clk_i as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7753__A1 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4567__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7748_ _3120_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7679_ _1385_ _1322_ _1394_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7808__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5819__A1 _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8481__A2 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__A2 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__C _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7441__B1 _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6795__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A2 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__A1 _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5030_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _3855_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7027__A3 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8224__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7060__I _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5038__A2 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6981_ _3907_ _1336_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7995__I _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7983__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6786__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7983__B2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5932_ _1392_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8720_ _0197_ clknet_leaf_77_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8651_ _0128_ clknet_leaf_75_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ _0461_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6538__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7735__A1 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7602_ _1177_ _3012_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_107_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4814_ _4095_ _0392_ _0403_ _0414_ _4060_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8582_ _0059_ clknet_leaf_67_wb_clk_i as2650.r123_2\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5794_ _1026_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7533_ _2942_ _2945_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _4189_ _4177_ _4172_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7464_ _2877_ _2878_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4676_ _4255_ _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8160__A1 _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8160__B2 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6415_ _1508_ _1861_ _1897_ _1762_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4859__I _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7395_ as2650.pc\[6\] _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6279__C _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput29 net53 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6346_ _1789_ _1798_ _1830_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4721__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6277_ _4234_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8016_ _2893_ _3363_ _3369_ _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5228_ _0797_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7018__A3 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5159_ _0739_ _0751_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5029__A2 _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7974__A1 _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__B2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7838__C _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8849_ net46 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8539__CLK clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4960__A1 _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8151__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7145__I _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6701__A2 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8454__A2 _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5268__A2 _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7662__B1 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5821__C _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8206__A2 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7965__A1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5440__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7717__A1 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _4097_ _4110_ _4017_ _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4951__A1 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4461_ as2650.addr_buff\[5\] _4041_ _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6200_ _1686_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7180_ _4224_ _4085_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4392_ _3972_ _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _1628_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8445__A2 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6456__A1 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7004__B _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _0533_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__I _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6759__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7956__A1 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7956__B2 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6223__A4 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6964_ _2376_ _2394_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8703_ _0180_ clknet_leaf_20_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5915_ _0587_ _0590_ _1432_ _0503_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7708__A1 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6895_ _0459_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6134__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5846_ _1031_ _1025_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8634_ _0111_ clknet_leaf_66_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7184__A2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8381__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ _4129_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8565_ _0042_ clknet_leaf_45_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6931__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7516_ _1317_ _2927_ _2929_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4728_ _4045_ _4222_ _0329_ _4042_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_124_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8496_ _2361_ _3821_ _3819_ _3822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8133__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7447_ _2521_ _2861_ _2862_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4659_ _4203_ _4209_ _4238_ _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6695__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7378_ _1332_ _2793_ _2794_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6329_ _0318_ _1812_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8436__A2 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6998__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7947__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8372__A1 _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7175__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8124__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4720__C _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__B _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4449__B1 _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6989__A2 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8704__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A1 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6219__I _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5110__B2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5661__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_29_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4962__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ _1111_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ _2137_ _2126_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5631_ _0741_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5177__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5793__I _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6913__A2 _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8350_ _3684_ _1472_ _3690_ _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5562_ as2650.stack\[1\]\[1\] _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8115__A1 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8102__C _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7301_ _0893_ _2717_ _2719_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4513_ _4093_ _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8281_ _2974_ _3623_ _3624_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5493_ as2650.pc\[1\] _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6677__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7232_ _2421_ _2638_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4444_ _4024_ _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7163_ _1081_ _1069_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4375_ _3954_ _3955_ _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6114_ _1024_ _1614_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7094_ _1377_ _2187_ _2513_ _2515_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6045_ _1546_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7669__B _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6573__B _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7996_ _3349_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _3958_ _3961_ _2377_ _2141_ _2263_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6878_ _2272_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8354__A1 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8617_ _0094_ clknet_leaf_56_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _1347_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4915__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8548_ _0025_ clknet_leaf_53_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5208__I _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8479_ _3806_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6668__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6132__A3 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8727__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8409__A2 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5891__A2 _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7093__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6039__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8345__A1 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7148__A2 _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8203__B _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4382__A2 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4957__I _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5331__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5882__A2 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7084__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5095__B1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6831__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4906__B _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4692__I _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7850_ _1112_ _3239_ _3244_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _0401_ _0547_ _0622_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5398__B2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4993_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7781_ _0865_ _2765_ _3182_ _3183_ _2286_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_90_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5937__A3 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6732_ _2184_ _1408_ _2153_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8336__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6663_ as2650.addr_buff\[1\] _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6347__B1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6898__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ as2650.stack\[2\]\[11\] _1170_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8402_ _2299_ _3733_ _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ as2650.r123_2\[0\]\[5\] _2044_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8333_ _3318_ _2156_ _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5570__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5545_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8264_ _2956_ _3609_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5476_ _1017_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4427_ _3969_ _4006_ _4007_ _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7215_ _2525_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8195_ _3541_ _3542_ _3454_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5873__A2 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7146_ _2554_ _2567_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4358_ _3902_ _3926_ _3938_ _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7077_ as2650.psu\[7\] _1641_ _2499_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4289_ _3869_ _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6822__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6028_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4535__C _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8007__C _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7979_ _3307_ _2600_ _3333_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8327__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout53 net29 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7418__I _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5313__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5313__B2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7066__A1 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6992__I _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5401__I _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_80 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_91 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6041__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8318__A1 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6232__I _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7541__A2 _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4355__A2 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ _0924_ as2650.stack\[3\]\[9\] as2650.stack\[2\]\[9\] _0908_ _0925_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4687__I _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _4131_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7000_ _2267_ _2425_ _2429_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5192_ _0657_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_44_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7057__A1 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__A2 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6280__A2 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7902_ as2650.stack\[3\]\[10\] _3275_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5311__I _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7833_ _3230_ _3232_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6032__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7764_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8309__A1 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4976_ _0476_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ net22 _2165_ _2168_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8572__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4594__A2 _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7695_ _1451_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6142__I _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6646_ _3898_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6577_ as2650.r123_2\[0\]\[2\] _2045_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8316_ _3559_ _3658_ _3659_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5528_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7296__A1 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8247_ net51 _3567_ _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5459_ _1043_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4649__A3 as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8178_ _3319_ _3511_ _3526_ _3167_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_59_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7048__A1 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7129_ _1051_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7599__A2 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7063__A4 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6271__A2 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4282__A1 _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7220__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6023__A2 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7771__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4424__I3 _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__A2 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5782__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6987__I _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8079__A3 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4300__I as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7039__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A4 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8251__A3 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_opt_2_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7767__B _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8595__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7211__A1 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _0428_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7486__C _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6565__A3 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7762__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5773__A1 _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _0362_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6500_ _1474_ _1761_ _1980_ _1705_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7480_ _2885_ _2887_ _2892_ _2894_ _2854_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_140_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4692_ _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7514__A2 _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6431_ _1848_ _1873_ _1894_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6362_ _1829_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5313_ _0905_ as2650.stack\[3\]\[8\] as2650.stack\[2\]\[8\] _0908_ _0909_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7278__A1 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8101_ _1509_ _3383_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6293_ _0816_ _4260_ _1733_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5244_ _0840_ _0826_ _0354_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8032_ _1513_ _3351_ _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8490__A3 _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _0739_ _0751_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7521__I _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6253__A2 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7450__A1 _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6005__A2 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7816_ _0855_ _3214_ _3216_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8796_ _0273_ clknet_3_1_0_wb_clk_i as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4567__A2 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7747_ _3131_ _0363_ _3149_ _3151_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5764__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4959_ _4161_ _0554_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7678_ _1502_ _2235_ _3084_ _3968_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_71_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7505__A2 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4319__A2 as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _1337_ _1400_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5819__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8481__A3 _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7441__A1 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7441__B2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6795__A3 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7992__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7587__B _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4790__I _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__B _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4730__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7680__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4494__A1 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__C _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7027__A4 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7432__A1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6980_ _2409_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6786__A3 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5931_ _1443_ _0830_ _1446_ _4229_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_111_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8650_ _0127_ clknet_leaf_72_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ _3967_ _3985_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7735__A2 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7601_ _1172_ _1165_ _2922_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_61_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4813_ _4078_ _0413_ _4094_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5746__A1 as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8581_ _0058_ clknet_leaf_62_wb_clk_i as2650.r123_2\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5793_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7532_ _2943_ _2944_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4744_ _0342_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7499__A1 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7463_ _2824_ _2830_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4675_ _4254_ _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8160__A2 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6414_ _0547_ _1861_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7394_ _2808_ _2810_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput19 net19 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6345_ _1793_ _1797_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4721__A2 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5036__I _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6276_ _1666_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8015_ _2608_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5227_ as2650.holding_reg\[7\] _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8760__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _0753_ _0754_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_57_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7423__A1 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ _0586_ _0539_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__A2 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4824__B _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8848_ net46 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8779_ _0256_ clknet_leaf_28_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8669__D _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8151__A2 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5268__A3 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7662__A1 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6465__A2 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7662__B2 _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7161__I _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4476__A1 _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4718__C _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7965__A2 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7717__A2 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8390__A2 _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ as2650.addr_buff\[6\] _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4391_ _3971_ _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6130_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6061_ _1574_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7653__A1 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6963_ _2216_ _2393_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8702_ _0179_ clknet_leaf_20_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5914_ _0678_ _0829_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6894_ _3975_ _2330_ _2334_ _2277_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_59_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7708__A2 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8633_ _0110_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5719__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5845_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8381__A2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6392__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8564_ _0041_ clknet_leaf_44_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5776_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7515_ _1634_ _2903_ _2928_ _2289_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_124_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4727_ _0326_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8495_ _3189_ _3102_ _1334_ _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8133__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7446_ _2812_ _2578_ _2579_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4658_ _4209_ _4237_ _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6695__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7377_ _0616_ _2089_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4589_ _4165_ _4168_ _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6328_ _4072_ _1665_ _1811_ _0307_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7644__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6259_ as2650.r0\[3\] _0525_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__A3 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7947__A2 _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5958__A1 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6325__I _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8656__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8372__A2 _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6060__I _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7635__A1 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6438__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7938__A2 _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5630_ _1163_ _1194_ _1196_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6374__A1 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5561_ _1137_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7300_ as2650.stack\[6\]\[3\] _2535_ _2718_ as2650.stack\[7\]\[3\] _2719_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6126__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4512_ _4076_ _3924_ _4058_ _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8280_ _3623_ _3624_ _2974_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5492_ _1067_ _1076_ _1079_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7231_ _2128_ _2473_ _2650_ _1323_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6677__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ as2650.psl\[3\] _4023_ _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4374_ net10 _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_119_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7162_ _1082_ _2582_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8529__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6113_ _1055_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7626__A1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7093_ _1035_ _1056_ _2280_ _2514_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5314__I _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6044_ _1368_ _1328_ _1545_ _1553_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8051__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8051__B2 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7995_ _3900_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6145__I _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _2101_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _3954_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5984__I _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8354__A2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8616_ _0093_ clknet_leaf_56_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5828_ _1059_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8547_ _0024_ clknet_leaf_59_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5759_ _1244_ _1275_ _1279_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4915__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6117__A1 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8478_ _2191_ _3801_ _3805_ _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6668__A2 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7429_ _2844_ _0534_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7704__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7093__A2 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8290__A1 _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6840__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7579__C _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4851__A1 _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8042__A1 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8345__A2 _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4504__S _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8203__C _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4303__I _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7856__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7608__A1 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7084__A2 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5095__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5095__B2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__A2 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6800_ _4234_ _0318_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_97_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6595__A1 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7780_ as2650.psu\[4\] _3111_ _3116_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4992_ _0587_ _0590_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5937__A4 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6731_ _2183_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8336__A2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6662_ _2071_ _2120_ _2124_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6347__A1 _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8401_ _3123_ _3732_ _3197_ _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _2057_ _2059_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5309__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8332_ _3343_ _3673_ _3674_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5544_ _1123_ _1125_ _1110_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5570__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8263_ _2474_ _3594_ _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5475_ _1023_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7524__I _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7214_ _2583_ _2634_ _2433_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4426_ as2650.holding_reg\[0\] _3980_ _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8194_ _1547_ _0803_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7145_ _2566_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4357_ _3927_ _3931_ _3937_ _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5044__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8272__A1 _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4288_ _3868_ _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7076_ _1641_ _1352_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6584__B _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5086__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6822__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6027_ _1534_ _1543_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_100_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__B1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7378__A3 _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6035__C2 _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7978_ _1511_ _2604_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4597__B1 _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6929_ _2353_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8304__B _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8327__A2 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8023__C _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7838__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7434__I _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7066__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8263__A1 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5077__A1 _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4793__I _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4824__A1 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6577__A1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_70 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_81 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_92 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6329__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5001__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7772__C _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5552__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4968__I _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7829__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5191_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8254__A1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5799__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6804__A2 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4815__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8006__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7901_ _3251_ _3273_ _3276_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7012__C _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7832_ _0870_ _2874_ _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6568__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7763_ _1414_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4975_ _0470_ _0473_ _0475_ _0476_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__8309__A2 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5240__A1 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6714_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5791__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7694_ _3098_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6645_ as2650.cycle\[7\] _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6740__A1 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6576_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8315_ net39 _3407_ _3614_ _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5527_ _1108_ _1109_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8246_ _3410_ _3591_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4409_ _3950_ _3979_ _3989_ _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8177_ _3366_ _3505_ _3525_ _2397_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ as2650.stack\[7\]\[13\] as2650.stack\[4\]\[13\] as2650.stack\[5\]\[13\] as2650.stack\[6\]\[13\]
+ _0884_ _0886_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7048__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7128_ _1069_ _2292_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5059__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7059_ _2373_ _2484_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5502__I _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A2 _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7220__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5231__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__A2 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8484__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7039__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8236__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6798__A1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7211__A2 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5222__A1 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7339__I _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _3998_ _0343_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5773__A2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _1848_ _1894_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6361_ _1831_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8100_ _1541_ _0557_ _3450_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_142_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8475__A1 _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6292_ _1727_ _1753_ _1777_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8031_ _1513_ _3351_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5243_ _0603_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8227__A1 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5174_ _0739_ _0751_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5322__I _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7450__A2 _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5461__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6581__C _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7202__A2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7815_ _0864_ _2821_ _3215_ _1493_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8795_ _0272_ clknet_3_1_0_wb_clk_i as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5213__A1 _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7746_ _3133_ _0337_ _3150_ _2474_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4958_ _4118_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5764__A2 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7677_ _2108_ _3083_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4889_ _0488_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6628_ _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6559_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8229_ _3512_ _3515_ _3575_ _3534_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8218__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7441__A2 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5452__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7587__C _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5204__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4638__S0 _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__B1 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4311__I as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8457__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7680__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4494__A2 _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7778__B _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5930_ _1432_ _1442_ _1445_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_81_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7069__I _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7196__A1 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7196__B2 _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8393__B1 _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7600_ _2612_ _2995_ _3008_ _2614_ _3010_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4812_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8580_ _0057_ clknet_3_5_0_wb_clk_i as2650.r123_2\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5792_ _1043_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ _2907_ _2913_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4743_ _4174_ _4181_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__S _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7462_ _2811_ _1489_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4674_ as2650.r123\[0\]\[1\] as2650.r123_2\[0\]\[1\] _3851_ _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6413_ _1806_ _1871_ _1872_ _1896_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7393_ _1116_ _2809_ _2191_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8448__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _1826_ _1827_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6275_ _1678_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7120__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8014_ _3319_ _3346_ _3367_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5226_ _4052_ _0822_ _4250_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5157_ _0625_ _4001_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5088_ _0357_ _0685_ _0358_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5434__A1 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8363__I _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7187__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8778_ _0255_ clknet_leaf_27_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5737__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7729_ _2492_ _4249_ _3134_ _3131_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7707__I _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__I as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8439__A1 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8585__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7111__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7442__I _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7662__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4476__A2 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6870__B1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6925__A1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5728__A2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4390_ _3970_ _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5900__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7653__A2 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input8_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ _0592_ _0608_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5416__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6962_ _2105_ _2383_ _2390_ _2392_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8701_ _0178_ clknet_leaf_26_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7020__C _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5913_ _0510_ _0610_ _0698_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6893_ _2139_ _2333_ _2330_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7169__A1 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8632_ _0109_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ _3933_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5719__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8563_ _0040_ clknet_leaf_44_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ _1289_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7514_ _2292_ _2914_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4726_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8494_ _3814_ _3819_ _3952_ _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7445_ _2523_ _2857_ _2860_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4657_ _4211_ _4223_ _4236_ _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7341__A1 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7376_ _3934_ _1051_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7892__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4588_ _3970_ _4166_ _4167_ _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6327_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6258_ _0742_ _1743_ _1744_ _0786_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5655__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5209_ net3 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _1666_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5407__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8093__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__A2 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5894__A1 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8268__I _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4796__I _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7172__I _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7635__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5646__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4449__A2 _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7399__A1 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4745__B _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7399__B2 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6071__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8600__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6374__A2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7571__A1 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _1076_ _1136_ _1139_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_38_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4511_ _4091_ _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7323__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5491_ as2650.stack\[0\]\[0\] _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6126__A2 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7230_ _0308_ _2599_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4442_ as2650.carry _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5885__A1 _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7161_ _2581_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4373_ _3953_ _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6112_ _1607_ _1609_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7626__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7092_ _1036_ _1038_ _1056_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _1555_ _1559_ _3848_ _1533_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_112_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7031__B _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7994_ _3322_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _2375_ _1612_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6876_ _2278_ _2298_ _2318_ _2277_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_74_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8615_ _0092_ clknet_leaf_53_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5827_ _0618_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__A1 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8546_ _0023_ clknet_leaf_57_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5758_ as2650.stack\[4\]\[6\] _1277_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6117__A2 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8477_ _0938_ _2636_ _3802_ _3804_ _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5689_ _1228_ _1230_ _1231_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7428_ _0615_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7359_ as2650.pc\[5\] net1 _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7078__B1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__A2 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8290__A2 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8623__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4565__B _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8037__B _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A2 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8042__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7250__B1 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8773__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4603__A2 _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5800__A1 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6356__A2 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7167__I _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4367__A1 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7305__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7856__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__I1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5867__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5619__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8281__A2 _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6044__A1 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4991_ as2650.holding_reg\[5\] _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7792__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6730_ _1026_ _3906_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_63_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8336__A3 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6661_ _2122_ _2123_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7544__A1 _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6347__A2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4358__A1 _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5612_ _1178_ _1179_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8400_ _1478_ _1473_ _2365_ _3731_ _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6910__S _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6592_ _0519_ _2032_ _2058_ _2054_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8331_ net40 _3407_ _3614_ _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8262_ _2915_ _2946_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7847__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5474_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5402__S0 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7213_ _2471_ _2584_ _2632_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7026__B _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ _4005_ _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8193_ _3539_ _3521_ _3540_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5325__I _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7144_ _2146_ _1616_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8646__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__A1 _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4356_ _3933_ _3936_ _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8272__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _1406_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4287_ as2650.ins_reg\[6\] _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6283__A1 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5086__A2 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7480__B1 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6026_ _1537_ _1540_ _1542_ _3847_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_74_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8796__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6035__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__B2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7977_ _2300_ _2615_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5995__I _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7783__A1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6928_ _2363_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ _1365_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6338__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__B _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8529_ _0006_ clknet_leaf_76_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5849__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8693__D _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5077__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__A1 _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_60 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__A2 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7774__A1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_71 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_82 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_93 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7526__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__I as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4760__A1 _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7829__A2 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6501__A2 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4512__A1 _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ as2650.r123\[0\]\[7\] as2650.r123_2\[0\]\[7\] _3851_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8456__I _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8254__A2 _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4815__A2 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7900_ as2650.stack\[3\]\[9\] _3275_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7831_ _1957_ _2286_ _1494_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6568__A2 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7765__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6704__I _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4579__A1 _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4974_ _0570_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7762_ _2323_ _0390_ _2436_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5240__A2 _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_53_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6713_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7693_ _3099_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _1363_ _4130_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8190__A1 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _0848_ _2005_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6740__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8314_ _1178_ _3409_ _3653_ _3657_ _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5526_ _1013_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4751__A1 _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8245_ _3365_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5457_ _4019_ _4102_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4503__A1 _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4408_ _3985_ _3988_ _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8176_ _3518_ _3524_ _2327_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5388_ _0649_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6595__B _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8366__I _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7127_ _2548_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4894__I _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7048__A3 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4339_ _3912_ _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5059__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7058_ as2650.cycle\[5\] _2483_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4806__A2 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _0817_ _1434_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6008__A1 _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7756__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7508__A1 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8181__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4742__A1 _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8484__A2 _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7039__A3 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8236__A2 _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4753__B _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7747__A1 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6524__I _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4690_ as2650.r0\[3\] _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7355__I _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6360_ _1836_ _1844_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4733__A1 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5311_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6291_ _1730_ _1752_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8475__A2 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8030_ _3977_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5242_ _4015_ _0833_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8227__A2 _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5173_ _0768_ _0755_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7986__A1 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5461__A2 _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4663__B _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7738__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7814_ _1197_ _3156_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8794_ _0271_ clknet_leaf_11_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7745_ _3133_ _0331_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5764__A3 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4972__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7676_ _3082_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4888_ _0486_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8163__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4889__I _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6627_ _1386_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7910__A1 as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _1606_ _0856_ _1652_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ _1094_ _1084_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6489_ _0816_ _1957_ _1921_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6477__A1 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8228_ _0806_ _0821_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7214__B _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8159_ _2832_ _3507_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6229__A1 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7977__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7729__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8045__B _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__S1 _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4963__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8154__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7901__A1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6947__C _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8707__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5691__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _1376_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7196__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8393__A1 _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8393__B2 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4811_ _0405_ _0407_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _1307_ _1309_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7530_ _2937_ _0714_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4954__A1 _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4742_ _4168_ _4172_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7461_ _1129_ _1550_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4673_ _4150_ _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6412_ _1719_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7392_ _2519_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6343_ _1782_ _1788_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6459__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6274_ _3901_ _1691_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7120__A2 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8013_ _3347_ _3362_ _3364_ _3366_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6429__I _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5225_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5156_ _0532_ _4255_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7959__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ _3974_ _0682_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_99_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6631__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5434__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7187__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8384__A1 _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8777_ _0254_ clknet_leaf_28_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _1470_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4945__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7728_ _3133_ _4245_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8136__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8312__C _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7659_ _3065_ _3066_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5508__I _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6698__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4412__I _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8439__A2 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5370__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6870__A1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5189__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8503__B _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6925__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8127__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4322__I _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _3998_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5664__A2 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7789__B _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__B1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6613__A1 as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5416__A2 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6961_ _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8700_ _0177_ clknet_leaf_26_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ _0456_ _1429_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6892_ _2144_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7169__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8631_ _0108_ clknet_leaf_12_wb_clk_i as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5843_ as2650.psl\[6\] _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6712__I _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8562_ _0039_ clknet_leaf_46_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8118__A1 _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5774_ _1286_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7513_ _2560_ _2926_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4725_ _4083_ _4086_ _4089_ _4006_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_8493_ _3818_ _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4656_ _4225_ _4228_ _4235_ _4074_ _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7444_ _2858_ _2859_ _2814_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5352__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__B2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ as2650.holding_reg\[1\] _3970_ _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7375_ _1115_ _2791_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6326_ _3948_ _1659_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5104__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6257_ _3999_ _0788_ _0744_ _0561_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6852__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5655__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _4070_ _1674_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5998__I _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ _0664_ _0735_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_131_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A2 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5958__A3 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6080__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8357__A1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6622__I _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8109__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8552__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7096__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5646__A2 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5701__I _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7571__A2 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _4090_ _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5490_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8520__A1 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5334__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4987__I as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ _4021_ _4020_ _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5885__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7160_ _2259_ _2506_ _2510_ _2518_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_119_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4372_ as2650.halted _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7087__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6111_ _1611_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7091_ _2512_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _0896_ _1556_ _1557_ _1558_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_140_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7993_ _2226_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6944_ _2170_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8339__A1 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6875_ _1609_ _2317_ _2298_ _2174_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7011__A1 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8614_ _0091_ clknet_leaf_53_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5826_ _0613_ _0460_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5022__B1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5573__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8545_ _0022_ clknet_leaf_56_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4376__A2 _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5757_ _1242_ _1275_ _1278_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4708_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8476_ _2620_ _2337_ _3803_ _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5688_ as2650.stack\[2\]\[0\] _1195_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8511__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7427_ _0712_ _0629_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _4087_ _4218_ _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7358_ _2572_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7078__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5007__B _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7078__B2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6309_ _1791_ _1794_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7289_ net8 _0296_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_77_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5521__I _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8042__A3 _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5800__A2 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7002__A1 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8502__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5316__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7183__I _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5867__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8266__B1 _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6816__A1 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7084__A4 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8018__B1 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8598__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7241__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6044__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7792__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7358__I _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6660_ _2118_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ _0472_ _1110_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4358__A2 _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6591_ _0973_ _2048_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8330_ _1185_ _3377_ _3672_ _2331_ _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5542_ _0710_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8261_ _2367_ _2458_ _3601_ _3606_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5473_ _1050_ _1060_ _3986_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4510__I _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4424_ _4000_ _4002_ _4003_ _4004_ _3843_ as2650.ins_reg\[1\] _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__5402__S1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7212_ _2520_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8192_ _1488_ _0708_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4355_ _3934_ _3935_ _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7143_ _2564_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4530__A2 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6807__A1 _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7074_ _2434_ _3928_ _2479_ _2497_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ _3866_ _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4666__B _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7480__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6283__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ as2650.psl\[1\] _4225_ _1541_ _3951_ _1484_ _1361_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__7480__B2 _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5341__I _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6035__A2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ _3321_ _3329_ _3330_ _3307_ _3167_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7783__A2 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6927_ _0485_ _2362_ _2353_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4597__A2 _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6858_ net25 _2300_ _2181_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ _1325_ _4143_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_52_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6789_ _2111_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8528_ _0005_ clknet_leaf_76_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8459_ _1018_ _0942_ _2424_ _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5516__I _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5849__A2 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7731__I _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7471__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8740__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5251__I _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7223__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_61 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_72 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_83 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A2 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_94 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__7178__I _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8511__B _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5426__I _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4760__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A2 _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7641__I _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7462__A1 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__B _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7830_ _1299_ _3114_ _3229_ _0856_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7765__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4579__A2 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7761_ _2492_ _0422_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4973_ _0470_ _0571_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6206__B _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6712_ _3955_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8309__A4 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7692_ _3098_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ _2102_ _2104_ _2105_ _1502_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_32_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8190__A2 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6574_ _2042_ _2043_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8313_ _3654_ _3656_ _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5525_ _0520_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4751__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8244_ _3559_ _3589_ _3590_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5456_ _3873_ _3867_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8794__D _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4407_ _3883_ _3987_ _3988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8763__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8175_ _3357_ _3522_ _3523_ _1708_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5387_ as2650.r123\[0\]\[5\] _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _2546_ _2547_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4338_ _3912_ _3887_ _3918_ _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_101_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6256__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7453__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7057_ _2480_ _2481_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4269_ as2650.halted net10 _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6008_ _3966_ _0844_ _1452_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7205__A1 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6008__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7205__B2 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7756__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7959_ _2220_ _2230_ _2506_ _3313_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7508__A2 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7726__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8469__B1 _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4742__A2 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7141__B1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6247__A2 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7444__A1 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6805__I _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7747__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6026__B _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8636__CLK clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A1 _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8786__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4733__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5310_ _0889_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6290_ _1774_ _1754_ _1775_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7683__A1 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ _4022_ _0835_ _0837_ _0351_ _4183_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_88_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5172_ _0612_ _4259_ _0753_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7435__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6916__S _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7986__A2 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7738__A2 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7813_ _3212_ _3138_ _3213_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5749__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8793_ _0270_ clknet_3_2_0_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7744_ _2107_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _0555_ _0514_ _0515_ _0378_ _0379_ _0499_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_33_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7675_ as2650.addr_buff\[7\] _3936_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4972__A2 _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _0446_ _0413_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8163__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6626_ _1034_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6174__A1 _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7910__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6557_ _2026_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5921__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _0949_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6488_ _1955_ _1962_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7674__A1 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8227_ _2552_ _3573_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_79_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5439_ _3881_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8158_ _3503_ _3506_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8218__A3 _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7426__A1 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6229__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ _0874_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8089_ _2686_ _3411_ _3439_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__A2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8326__B _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8659__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4660__A1 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7729__A2 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6401__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8154__A2 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7201__I1 as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7901__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5912__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6468__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7665__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7191__I _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5704__I _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7417__A1 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8236__B _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4651__A1 _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8393__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4810_ _0410_ _3860_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _1308_ _1284_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4403__A1 _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4954__A2 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7460_ _2528_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4672_ _4162_ _4195_ _4251_ _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ _1848_ _1875_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_70_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5903__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7391_ _2772_ _2807_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6342_ _1782_ _1788_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6459__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6273_ _1692_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8012_ _3365_ _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5224_ _0797_ _0379_ _0798_ _0555_ _0801_ _0378_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_102_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5155_ _0563_ _0747_ _0752_ _0660_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_69_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7959__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8081__A1 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8801__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5086_ _0683_ _0443_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8146__B _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7050__B _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6631__A2 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8384__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8776_ _0253_ clknet_leaf_27_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6395__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _1485_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7727_ _2401_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4939_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4945__A2 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8136__A2 _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6180__I _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7658_ as2650.pc\[13\] _1184_ _2993_ _2994_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _3895_ _3881_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6698__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7589_ as2650.addr_buff\[3\] _2998_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_opt_1_0_wb_clk_i clknet_3_3_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8439__A3 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5370__A2 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7647__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8072__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8375__A2 _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8127__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7914__I _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4759__B _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7638__A1 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6974__B _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6466__S _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4872__B2 _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8063__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7810__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6960_ _2179_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _4037_ _4195_ _0363_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_59_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ _3976_ _2330_ _2332_ _2277_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7169__A3 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8630_ _0107_ clknet_leaf_12_wb_clk_i as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5842_ _1358_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8561_ _0038_ clknet_leaf_49_wb_clk_i as2650.stack\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5773_ _3884_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8118__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7512_ _2122_ _2380_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6129__A1 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4724_ _0309_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8492_ _1310_ _3815_ _3816_ _3817_ _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7443_ _2822_ _2833_ _2775_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4655_ _4227_ _4234_ _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7374_ _2730_ _2741_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ _4083_ _4086_ _4089_ _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_116_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7629__A1 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6325_ _1686_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5344__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6256_ as2650.r0\[1\] _0787_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6301__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _0635_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6852__A2 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6187_ _1365_ _1385_ _1672_ _1673_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_69_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8054__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5138_ _0667_ _0668_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6175__I _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7801__A1 _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5069_ _0409_ _4255_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8323__C _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8759_ _0236_ clknet_leaf_42_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5040__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7096__A2 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8293__A1 _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8293__B2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4854__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8045__A1 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8348__A2 _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6813__I _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6359__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5031__A1 _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6969__B _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8520__A2 _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4440_ _3982_ _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6531__A1 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5334__A2 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ _3951_ _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6110_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8284__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7090_ _3910_ _1326_ _2241_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5098__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ as2650.psu\[4\] _1541_ _1484_ net27 _0883_ _1539_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8036__A1 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7992_ _3345_ _2597_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_96_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6943_ _2163_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4952__B _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5270__A1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6723__I _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6874_ _2299_ _2314_ _2315_ _2316_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4671__C _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7011__A2 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8613_ _0090_ clknet_leaf_52_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5825_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5022__A1 _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8544_ _0021_ clknet_leaf_56_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5756_ as2650.stack\[4\]\[5\] _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5573__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4707_ _4215_ _4217_ _4219_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8475_ _3795_ _2336_ _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5687_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8511__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7426_ _2811_ _2841_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4638_ as2650.r123\[1\]\[2\] as2650.r123\[0\]\[2\] as2650.r123_2\[1\]\[2\] as2650.r123_2\[0\]\[2\]
+ _3843_ _3853_ _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6522__A1 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7357_ _1115_ _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_85_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4569_ _4128_ _4136_ _4149_ _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8275__A1 _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7078__A2 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _0292_ _0744_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7288_ _0304_ _4216_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5089__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8385__I as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6239_ _0627_ _4259_ _0776_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4836__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8027__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6038__B1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6589__A1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7250__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8334__B _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5261__A1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5800__A3 _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7002__A2 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5564__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__A3 _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6513__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7710__B1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8266__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8509__B _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8018__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8018__B2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4328__I _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7241__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6201__B1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5610_ _1084_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6590_ _1908_ _2028_ _2034_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4358__A3 _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ as2650.pc\[6\] _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8260_ _3603_ _3605_ _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5472_ _0357_ _1051_ _1057_ _1058_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7211_ _2594_ _2619_ _2631_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4423_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] _3852_ _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8191_ _1488_ _0708_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8257__A1 _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7142_ _0459_ _1611_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4354_ as2650.addr_buff\[6\] _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6807__A2 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7073_ _3885_ _2458_ _2494_ _2496_ _2164_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4285_ as2650.ins_reg\[4\] _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_140_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8009__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _0542_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__A2 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7975_ _2233_ _2226_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _2133_ _2360_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _2083_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5808_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6788_ _1369_ _1380_ _1308_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5546__A2 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8527_ _0004_ clknet_leaf_75_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5739_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4701__I _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8458_ _0937_ _1295_ _2352_ _3787_ _2593_ _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7409_ _1114_ net1 _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5849__A3 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8389_ _1333_ _1328_ _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8248__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5532__I _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7471__A2 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7223__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6026__A3 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5234__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_62 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_73 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_84 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6734__A1 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7194__I _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5707__I _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8487__A1 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8487__B2 _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8239__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A3 _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8565__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7462__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6273__I _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7760_ _2437_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4972_ _0409_ _4001_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6973__A1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _2164_ _1410_ _1319_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_75_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7691_ _1397_ _3079_ _3081_ _3097_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_71_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6642_ _1311_ _1616_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6725__A1 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _4198_ _2033_ _2030_ _0928_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8312_ _1178_ _3495_ _3497_ _3655_ _2320_ _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8478__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8243_ net51 _3557_ _3472_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5455_ _3940_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7150__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6876__C _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_62_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4406_ _3986_ _3862_ _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8174_ _1489_ _3083_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5386_ _0966_ _0860_ _0976_ _0977_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ _0459_ _2247_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4337_ _3914_ _3917_ _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7056_ _2480_ _2481_ _2482_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4268_ _3848_ _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6007_ _1360_ _1427_ _1524_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8402__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5216__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6183__I _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6964__A1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7958_ _3964_ _2116_ _2187_ _2232_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__5767__A2 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _2345_ _2347_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7889_ _3256_ _3264_ _3269_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5519__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__A1 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8469__A1 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8588__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7141__A1 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7141__B2 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8522__B _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6707__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6042__B _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5930__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7132__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ _0595_ _4109_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _0612_ _4259_ _0753_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7435__A2 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5446__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4516__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7812_ _1361_ _3110_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8792_ _0269_ clknet_leaf_16_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5749__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ _1086_ _3130_ _3136_ _3148_ _2372_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4955_ _0377_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_80_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__I _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7674_ _3080_ _1607_ _4049_ _2114_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_32_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ _0485_ _0461_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ _2080_ _2082_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_123_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5347__I _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7371__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ _2026_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5507_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6487_ _1952_ _1964_ _1967_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8226_ _3570_ _3572_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5438_ _3895_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7674__A2 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8157_ _2385_ _3505_ _2837_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5369_ _0391_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7108_ _0891_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7426__A2 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8088_ _2683_ _0393_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7039_ _2413_ _2154_ _2464_ _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_60_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8139__B1 _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7737__I _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7665__A2 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7417__A2 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5428__A1 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__I _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8603__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4651__A2 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8753__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _0340_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4671_ _4241_ _4246_ _4249_ _4052_ _4250_ _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7353__A1 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ _1890_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7390_ _2774_ _2783_ _2806_ _2727_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5903__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _1787_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6500__B _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ _1704_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8011_ _2233_ _2077_ _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5223_ _4201_ _0803_ _0819_ _4119_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6927__S _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5154_ _4213_ _0562_ _0567_ _0561_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6726__I _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8081__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5085_ as2650.holding_reg\[6\] _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7985__C _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8775_ _0252_ clknet_leaf_28_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7592__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ _0808_ _1501_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7726_ _2107_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4938_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4869_ _4080_ _3999_ _0367_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7344__A1 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7657_ as2650.pc\[14\] _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6608_ _1539_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6698__A3 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7588_ _2131_ _2998_ _2175_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7895__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7506__B _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6539_ _2007_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5805__I _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5107__B1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7647__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5658__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8209_ _3316_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8626__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8072__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8776__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7583__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4397__A1 _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7335__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7886__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5897__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5715__I _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6974__C _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A1 _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4872__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8063__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4494__C _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6074__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ _0831_ _0843_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6890_ _2137_ _2331_ _2330_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5841_ _1281_ _1341_ _1356_ _1359_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7574__A1 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5772_ _1288_ _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8560_ _0037_ clknet_leaf_49_wb_clk_i as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7511_ _2922_ _2924_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4723_ _4044_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8491_ _1297_ _1348_ _2498_ _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6129__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7326__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7442_ _2320_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4654_ _4185_ _4233_ _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5888__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7373_ _2785_ _2786_ _2788_ _2789_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_4585_ _4163_ _4164_ _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8649__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6324_ _1696_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4560__A1 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6255_ _1739_ _1741_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6301__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5104__A3 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4312__A1 _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5206_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6186_ _1659_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8799__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4863__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8054__A2 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5137_ _0667_ _0668_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5068_ _0665_ _0659_ _0666_ _0564_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5812__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4379__A1 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4704__I _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8758_ _0235_ clknet_leaf_43_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5040__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _0864_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7317__A1 _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8689_ _0166_ clknet_leaf_10_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5963__C _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5879__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8067__B _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6056__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8514__C _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__A1 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5031__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6969__C _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7859__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6531__A2 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _3856_ _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5098__A2 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ as2650.psu\[7\] _0807_ _1535_ as2650.psu\[5\] _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6276__I _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6047__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7991_ as2650.pc\[0\] _4063_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6598__A2 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7795__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6942_ _2373_ _2218_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5270__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_16_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6873_ _2107_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8612_ _0089_ clknet_leaf_52_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7011__A3 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5824_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5022__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8543_ _0020_ clknet_leaf_56_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5755_ _1268_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5686_ _1153_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8474_ _3783_ _3800_ _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7425_ _1114_ _1106_ _2741_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4637_ _4084_ _4216_ _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5355__I _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6522__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4533__A1 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7356_ _1107_ _1099_ _2684_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4568_ _3848_ _4148_ _4149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _1746_ _1790_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8275__A2 _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7287_ _2444_ _2685_ _2705_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4499_ _4079_ _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5089__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6238_ _1723_ _1724_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7483__B1 _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7503__C _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6186__I _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6169_ _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6038__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6038__B2 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5261__A2 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7538__A1 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4434__I _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6761__A2 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6513__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7710__A1 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8266__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6096__I _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8018__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7777__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7529__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6201__A1 _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6752__A2 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5540_ _1105_ _1120_ _1122_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ _3884_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7701__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ as2650.r123\[1\]\[0\] as2650.r123_2\[1\]\[0\] _3852_ _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4515__A1 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7210_ _2620_ _2584_ _2629_ _2630_ _2320_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8190_ _2305_ _3350_ _3323_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7604__B _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7141_ _2549_ _2550_ _2562_ _2344_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8257__A2 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4353_ as2650.addr_buff\[5\] _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7072_ _3928_ _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4284_ _3864_ _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _1538_ _0807_ _1539_ _4023_ as2650.overflow _0307_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__8009__A2 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7768__B2 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7974_ _3323_ _3325_ _3328_ _2485_ _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_81_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6925_ _0519_ _1527_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7766__S _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6856_ _1503_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5807_ _3920_ _3940_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6787_ _2031_ _1608_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7940__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8526_ _0003_ clknet_leaf_75_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4754__A1 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5738_ _1011_ _1151_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4754__B2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8457_ _1352_ _2350_ _1295_ _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5669_ as2650.r123_2\[3\]\[0\] _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4506__A1 _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7408_ _2823_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8388_ _1378_ _2229_ _3719_ _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7339_ _2530_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5813__I _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6259__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7208__B1 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7759__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8345__B _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5234__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_63 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_74 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_85 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6982__A2 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8080__B _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A1 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8487__A2 _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6819__I _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8239__A2 _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7998__A1 _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__B _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4681__B1 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _0293_ _4254_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6710_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7690_ _3085_ _3087_ _3093_ _3096_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_32_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6641_ _1392_ _2103_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6725__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4736__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6572_ as2650.r123_2\[0\]\[1\] _2027_ _2040_ _2041_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8311_ _2436_ _3646_ _3009_ _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5523_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6489__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _1035_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8242_ _2937_ _3344_ _3584_ _3374_ _3588_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_117_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7150__A2 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _3850_ _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8173_ _0714_ _0709_ _3521_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5385_ _0849_ _4148_ _0560_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7124_ _2085_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4336_ _3868_ _3916_ _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7055_ _2480_ _2481_ _2168_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4267_ _3847_ _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6661__A1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6006_ _1454_ _1466_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6413__A1 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5216__A2 _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7957_ _0460_ _2306_ _3311_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4975__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6908_ _4197_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7888_ as2650.stack\[4\]\[11\] _3266_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ _1033_ _2084_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5808__I _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4712__I _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7228__C _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8509_ _1286_ _3771_ _2346_ _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8469__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5527__I0 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7141__A2 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6639__I _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7244__B _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5543__I _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6955__A2 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8157__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6707__A2 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__I _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7380__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8532__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7132__A2 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7683__A3 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8682__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5170_ _0731_ _0757_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6993__B _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6643__A1 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8396__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7811_ net27 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8791_ _0268_ clknet_leaf_16_wb_clk_i net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7742_ _1472_ _3137_ _3147_ _2159_ _3098_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_127_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8148__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4954_ _4040_ _0518_ _0553_ _0334_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8148__B2 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7673_ _2097_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ as2650.holding_reg\[4\] _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6624_ _3962_ _2086_ _3955_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5382__A1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _0848_ _2005_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6887__C _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5506_ as2650.pc\[2\] _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8320__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6486_ _1953_ _1963_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8225_ _3082_ _3571_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5437_ _3906_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7674__A3 _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6882__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8156_ net34 _3504_ _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5368_ _0918_ _0956_ _0958_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7107_ _2528_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4319_ as2650.idx_ctrl\[1\] as2650.idx_ctrl\[0\] _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8087_ _3408_ _3437_ _3438_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5299_ _0874_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7038_ _2305_ _3984_ _2465_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8387__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6937__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8139__A1 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8139__B2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8311__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5125__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7417__A3 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5428__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6625__A1 _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8378__A1 _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7050__A1 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6832__I _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5448__I _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4352__I _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ _4138_ _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5364__A1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5364__B2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6340_ _1783_ _1800_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8302__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6500__C _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6271_ _1701_ _1713_ _1718_ _1757_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6864__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8010_ _2409_ _3363_ _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5667__A2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5222_ _4061_ _0815_ _0818_ _4201_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5153_ _0746_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7612__B _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6616__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5084_ _0676_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6092__A2 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8369__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8443__B _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7041__A1 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6742__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8774_ _0251_ clknet_leaf_27_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7592__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7725_ _2850_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4937_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7656_ _3063_ _3064_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4868_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _2068_ _0967_ _2040_ _2070_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7587_ _2919_ _2890_ _2997_ _2152_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ _4205_ _0312_ _0328_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6538_ _1822_ _2002_ _2013_ _2014_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6189__I _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5107__A1 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__B2 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6469_ _1916_ _1936_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6855__A1 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8208_ _2864_ _3344_ _3551_ _3374_ _3555_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5658__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8139_ _3378_ _3475_ _3488_ _3347_ _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6607__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8072__A3 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7280__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7748__I _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7032__A1 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5043__B1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7583__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4397__A2 _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7335__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__A2 _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__B _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6099__I _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5649__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4321__A2 _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8720__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7023__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5840_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7574__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4388__A2 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _3945_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7510_ _1159_ _2923_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _4220_ _0313_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8490_ _2163_ _1607_ _3721_ _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_124_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7326__A2 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5337__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7441_ _2636_ _2814_ _2821_ _2529_ _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6534__B1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ _4231_ _4232_ _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5888__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7372_ as2650.stack\[6\]\[5\] _2540_ _2718_ as2650.stack\[7\]\[5\] _0880_ _2789_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4584_ _3996_ _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6323_ _1807_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4560__A2 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6837__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _1731_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_103_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _0797_ _0419_ _0798_ _0512_ _0801_ _0418_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_131_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _1313_ _1335_ _3904_ _1032_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_69_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _0655_ _0730_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7262__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ _4080_ _0469_ _0567_ _0657_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7565__A2 _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8757_ _0234_ clknet_leaf_52_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5969_ _0711_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7708_ _0885_ _3114_ _2038_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8688_ _0165_ clknet_leaf_10_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8514__A1 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8514__B2 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5328__A1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7639_ _2935_ _3046_ _3048_ _2520_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5816__I _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5879__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__B _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__A2 _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5500__A1 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6056__A2 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8450__B1 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7253__B2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7478__I _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7800__I0 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5567__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8505__A1 _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6331__B _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6531__A3 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4542__A2 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8258__B _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6047__A2 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7990_ _3318_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7795__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _2372_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6872_ _1041_ _2307_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_50_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8611_ _0088_ clknet_leaf_52_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5823_ _1052_ _3933_ _4164_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8542_ _0019_ clknet_leaf_57_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_56_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5754_ _1239_ _1275_ _1276_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8616__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4705_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6507__B1 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8473_ _3786_ _3800_ _0943_ _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5685_ _1075_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8012__I _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7424_ _2612_ _2814_ _2835_ _2839_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4636_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _3853_ _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8766__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7355_ _2581_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4567_ _4138_ _4147_ _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6306_ _0785_ _1791_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8275__A3 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7286_ _2614_ _2692_ _2704_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8168__B _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4498_ as2650.r0\[1\] _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6286__A2 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7483__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _0770_ _0794_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7483__B2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4297__A1 _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6168_ _1654_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6038__A2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _0715_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _1593_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5320__B _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_57_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7710__A2 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8078__B _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7474__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6377__I _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7226__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7777__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A1 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6201__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5470_ _1008_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7701__A2 _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4421_ _4001_ _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4515__A2 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7671__I _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7140_ _2417_ _2556_ _2561_ _2086_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7604__C _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4352_ _3932_ _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7465__A1 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7071_ _2075_ _2488_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5191__I _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4283_ _3863_ _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6022_ _4064_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7217__A1 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7768__A2 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8435__C _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7973_ _2071_ _3327_ _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5779__A1 as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6976__B1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6924_ _1532_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _2248_ _2297_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8193__A2 _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5806_ _3983_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6786_ _1083_ _1309_ _2229_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7940__A2 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7067__B _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8525_ _0002_ clknet_leaf_72_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5737_ _1023_ _1061_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5951__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8456_ _3783_ _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5668_ _1138_ _1200_ _1219_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7407_ as2650.pc\[6\] net2 _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4506__A2 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _3989_ _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5703__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8387_ _0351_ _2091_ _2216_ _1388_ _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5599_ _1154_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7338_ _2549_ _2742_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6259__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7456__A1 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6197__I _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7269_ _2686_ _2687_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5050__B _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_64 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_75 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_86 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__I _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6195__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7931__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5942__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__I as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4745__A2 _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_1_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7491__I _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7424__C _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7447__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7998__A2 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6835__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4681__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8255__C _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4681__B2 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _0563_ _0564_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4433__A1 _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8702__D _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _1047_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7922__A2 _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6571_ _1771_ _2026_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4736__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8310_ _2915_ _3008_ _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5522_ as2650.pc\[4\] _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8241_ _2522_ _3587_ _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6489__A2 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5453_ _1036_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4404_ _3943_ _3981_ _3984_ _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7334__C _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8172_ _3519_ _3484_ _3520_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5384_ _0933_ _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7123_ _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4335_ _3915_ _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_87_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7054_ _2163_ _3891_ _1037_ _1028_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_59_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4266_ _3846_ _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6005_ _1500_ _1505_ _1522_ _1426_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6661__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4672__A1 _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6413__A2 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4265__I _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7610__A1 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7956_ _4140_ _3309_ _3310_ _2216_ _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_71_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _1482_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7887_ _3254_ _3264_ _3268_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _1032_ _3882_ _3960_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6177__A1 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5924__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6769_ _0466_ _1990_ _2213_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8508_ _3828_ _3830_ _3831_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7677__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7525__B _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8439_ _2272_ _2294_ _2511_ _3768_ _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_104_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5527__I1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7244__C _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5045__B _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6101__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__B _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4663__A1 _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7601__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8157__A2 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4903__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7904__A2 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__A2 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5915__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7668__A1 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6891__A2 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6993__C _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7840__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4654__A1 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 io_in[5] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7810_ _3132_ _3208_ _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8790_ _0267_ clknet_leaf_16_wb_clk_i net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4406__A1 _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _2448_ _1763_ _3146_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4953_ _0520_ _4062_ _0551_ _0552_ _4039_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7396__I _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8148__A2 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7672_ _3870_ _1450_ _4082_ _2279_ _3078_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4884_ _4160_ _0457_ _0484_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6623_ _2083_ _2085_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5906__A1 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _1999_ _2002_ _2025_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5382__A2 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5505_ _1067_ _1089_ _1091_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6485_ _1806_ _1949_ _1950_ _1966_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8020__I _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8224_ _1546_ _0802_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5436_ _3920_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6331__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7674__A4 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8155_ net52 _3474_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6882__A2 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5367_ _0910_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8084__A1 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7106_ _2179_ _1343_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4318_ _3889_ _3898_ _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8086_ net31 _3317_ _2938_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8176__B _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5298_ _0893_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7080__B _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ _2078_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7831__A1 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8387__A2 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4924__S _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7939_ _3282_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8139__A2 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7898__A1 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8311__A2 _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6322__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5125__A2 _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4884__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7702__C _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8086__B _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6625__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7822__A1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5222__C _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8378__A2 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7050__A2 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6334__B _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4633__I _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7889__A1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__A1 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5464__I _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6270_ _1719_ _1756_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _0817_ _4061_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6864__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4875__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8066__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5152_ _0747_ _0748_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6616__A2 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7813__A1 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5083_ _0678_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_96_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8443__C _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8773_ _0250_ clknet_leaf_27_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5985_ _1502_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4543__I _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8015__I _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7724_ _3101_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4936_ _0531_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_75_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7655_ _1191_ _2809_ _2168_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4867_ as2650.r123\[0\]\[3\] as2650.r123_2\[0\]\[3\] _0365_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6927__I0 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6606_ _1998_ _2045_ _2040_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7586_ as2650.addr_buff\[0\] as2650.addr_buff\[1\] as2650.addr_buff\[2\] _2997_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6552__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ _0316_ _0311_ _0314_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6537_ _0375_ _1912_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5374__I as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6304__A1 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5107__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ as2650.r123_2\[2\]\[5\] _1910_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8207_ _2732_ _2880_ _3554_ _2574_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7803__B _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5419_ _3883_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6399_ _0533_ _0741_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4866__A1 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8138_ _3481_ _3487_ _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6419__B _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6607__A2 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7804__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8069_ _0325_ _0330_ _0306_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_102_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7280__A2 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6933__I _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7032__A2 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5043__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5043__B2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8672__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4397__A3 _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7764__I _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6543__A1 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5284__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8048__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5282__A1 as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7939__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6843__I _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7023__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _3912_ _0850_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6999__B _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _0290_ _4199_ _4200_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7440_ _2822_ _2833_ _2840_ _2855_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5337__A2 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4652_ _3922_ _4068_ _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7371_ _0892_ _2787_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_122_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ _3994_ _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8287__A1 _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ _0464_ _1653_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4560__A3 _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6837__A2 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ as2650.r0\[5\] _0468_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4848__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _0797_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4848__B2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8039__A1 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7342__C _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6184_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8545__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5135_ _0656_ _0731_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4538__I _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7798__B1 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5066_ _0657_ _0471_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5812__A3 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8695__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5025__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5369__I _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4273__I _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6773__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8756_ _0233_ clknet_leaf_50_wb_clk_i as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5968_ _0847_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ _0410_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7707_ _3113_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5899_ _1414_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8687_ _0164_ clknet_leaf_10_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6525__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7638_ _2858_ _3047_ _3033_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7569_ _1316_ _2980_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8278__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4839__A1 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8450__A1 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8450__B2 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8202__A1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__I as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7708__B _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__I _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8505__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6516__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8269__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8568__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7443__B _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8441__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__A3 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5255__A1 _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6940_ _1357_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6871_ _2313_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5007__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5822_ _1293_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8610_ _0087_ clknet_leaf_11_wb_clk_i as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8541_ _0018_ clknet_leaf_53_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5753_ as2650.stack\[4\]\[4\] _1271_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4821__I _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__A1 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8472_ _1622_ _3766_ _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5684_ _1227_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6507__B2 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7423_ _2175_ _2838_ _2701_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4635_ _4214_ _3859_ _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7354_ _2373_ _2771_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_25_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _4139_ _4146_ _3989_ _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6305_ _4212_ _0788_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7285_ _1333_ _2702_ _2703_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4497_ _4077_ _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6236_ _0773_ _0793_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7483__A2 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4268__I _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6167_ _0464_ _1653_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _3923_ _0589_ _0619_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8432__A1 _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _1189_ _1600_ _1601_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5049_ _0638_ _0644_ _0647_ _3993_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6416__C _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8739_ _0216_ clknet_leaf_44_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5827__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8499__A1 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__A2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6658__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8078__C _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7474__A2 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5237__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6985__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5788__A2 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4641__I _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7162__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7952__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ as2650.r123\[0\]\[0\] as2650.r123_2\[0\]\[0\] _3852_ _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5712__A2 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7173__B _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _3887_ _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7070_ _2356_ _2492_ _2493_ _2464_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4282_ _3850_ _3862_ _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6021_ as2650.psl\[7\] _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7217__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__B _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6976__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7972_ _4047_ _3326_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5779__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6976__B2 _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6923_ _2359_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _2285_ _2287_ _2296_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6728__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_126_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5805_ _1053_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6785_ _4134_ _1409_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8524_ _0001_ clknet_leaf_72_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5736_ _1246_ _1258_ _1263_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5667_ as2650.stack\[1\]\[14\] _1135_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8455_ _1018_ _3784_ _3785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7153__A1 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _4197_ _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7406_ _3885_ _2814_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8386_ _1464_ _1451_ _1318_ _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6900__A1 _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5598_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5703__A2 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8179__B _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7083__B _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7337_ _2616_ _2750_ _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4549_ _4129_ _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7268_ as2650.pc\[3\] net8 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5315__C _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5467__A1 _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6219_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7199_ _2526_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8405__A1 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7102__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_54 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_65 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_76 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6941__I _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_87 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6719__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7258__B _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5557__I _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6195__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5942__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4902__B1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8606__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4681__A2 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6056__C _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8756__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__A2 _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7168__B _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7383__A1 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4371__I _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ _2039_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5521_ _1066_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7135__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8240_ _1159_ _3502_ _3586_ _2595_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5452_ _1027_ _1039_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4403_ _3982_ _3983_ _3915_ _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8171_ _2844_ _0642_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5383_ _0967_ _0973_ _0974_ _0951_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7122_ _2533_ _2537_ _2543_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4334_ as2650.ins_reg\[7\] _3915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ as2650.cycle\[4\] _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4265_ _3845_ _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6004_ _1506_ _1507_ _1510_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_45_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4672__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7955_ _3962_ _2086_ _2095_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6906_ _1628_ _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7886_ as2650.stack\[4\]\[10\] _3266_ _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6837_ _1025_ _2279_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7374__A1 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6177__A2 _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6768_ _0845_ _2195_ _2197_ as2650.r123\[2\]\[7\] _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7806__B _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8507_ _1443_ _3828_ _2167_ _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7126__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5719_ _1228_ _1250_ _1253_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6699_ _3958_ _4056_ _1039_ _1327_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8323__B1 _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8438_ _2514_ _3668_ _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7677__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8369_ _1117_ _3701_ _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6001__I _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8629__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7429__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6101__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6652__A3 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8779__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5860__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4663__A2 _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7601__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5612__A1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6671__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5287__I as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7365__A1 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5915__A2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7117__A1 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7668__A2 _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7007__I _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6846__I _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6643__A3 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7840__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5851__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 io_in[6] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4406__A2 _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4952_ _4095_ _0303_ _4060_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7740_ _1628_ _2176_ _3145_ _2424_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7671_ _2222_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4883_ as2650.r123\[1\]\[3\] _4151_ _0483_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _2084_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5906__A2 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4965__I0 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ as2650.r123_2\[1\]\[7\] _2015_ _2024_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5504_ as2650.stack\[0\]\[1\] _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6484_ _1912_ _1965_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7345__C _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7659__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8223_ _3539_ _3521_ _3569_ _3540_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5435_ _1018_ _1012_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6331__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8154_ _2160_ _2249_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5366_ _0905_ as2650.stack\[3\]\[11\] as2650.stack\[2\]\[11\] _0908_ _0959_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8457__B _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4317_ _3890_ _3894_ _3897_ _3898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7105_ _2526_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8085_ _2698_ _3409_ _3436_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5297_ _0892_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6095__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ _2325_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5142__I0 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7831__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7938_ _1232_ _3298_ _3299_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7869_ as2650.stack\[5\]\[11\] _3252_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7898__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6322__A2 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4884__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5833__A1 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7586__A1 as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5011__S _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6334__C _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A2 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7338__A1 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7889__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7446__B _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6561__A2 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8121__I _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7510__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5220_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4875__A2 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5151_ _0292_ _0562_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8066__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5480__I as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6077__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5082_ _0591_ _0599_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7813__A2 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7577__A1 _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8772_ _0249_ clknet_leaf_26_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _1376_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7723_ _1072_ _3100_ _3128_ _3129_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4935_ _0533_ _3860_ _4101_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7329__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7654_ _2471_ _3061_ _3062_ _3053_ _2682_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4866_ _4258_ _0374_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6927__I1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6605_ as2650.r123_2\[0\]\[7\] _2026_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6552__A2 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ _0382_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7585_ _2995_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4563__A1 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6536_ as2650.r123_2\[1\]\[2\] _2008_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6467_ _1808_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8206_ _2864_ _3502_ _3497_ _3553_ _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5418_ _1002_ _0860_ _1006_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6398_ _1880_ _1881_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5604__B _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8137_ _2136_ _3391_ _3486_ _2402_ _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5349_ _0900_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6607__A3 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7804__A2 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8068_ _3354_ _3418_ _3419_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5815__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7019_ _2426_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7568__A1 _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6543__A2 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7740__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8048__A2 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7256__B1 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4609__A2 _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7559__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4644__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _0291_ _4209_ _0321_ _4199_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _4068_ _4230_ _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5337__A3 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4582_ _4161_ _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7370_ _0898_ as2650.stack\[5\]\[5\] as2650.stack\[4\]\[5\] _2625_ _2787_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6321_ _1712_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6252_ as2650.r0\[6\] _0368_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5203_ _0634_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6183_ _1669_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8039__A2 _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5134_ _0663_ _0669_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7798__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7798__B2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5065_ _0532_ _4002_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6470__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4554__I _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8211__A2 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__A2 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6222__A1 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8755_ _0232_ clknet_leaf_50_wb_clk_i as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6773__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7970__A1 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7706_ _3846_ _1479_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4918_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8686_ _0163_ clknet_3_2_0_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_90_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5898_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7086__B _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7637_ _2768_ _3031_ _3034_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_138_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ _4180_ _0439_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4536__A1 _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7568_ _2663_ _2979_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6519_ _1808_ _1998_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8278__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7499_ _2909_ _2911_ _2912_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4839__A2 _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7105__I _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7789__A1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6944__I _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8450__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6461__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8202__A2 _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A1 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4775__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6516__A2 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8269__A2 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5244__B _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__I _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8441__A2 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__A4 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5255__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4374__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6870_ _1394_ _2301_ _2304_ _2312_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5007__A2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ _1295_ _1306_ _1331_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_35_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6755__A2 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8721__D _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8540_ _0017_ clknet_leaf_57_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5752_ _1266_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4703_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8471_ _3794_ _3799_ _2992_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5683_ as2650.r123_2\[3\]\[7\] _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6507__A2 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7422_ _2836_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4634_ _4213_ _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7180__A2 _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4565_ _4141_ _4142_ _4145_ _3862_ _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7353_ _2730_ _2582_ _2770_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5933__I _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7468__B1 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6304_ _1743_ _1747_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7284_ _0397_ _2101_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4496_ _4076_ _3919_ _4058_ _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6235_ _0765_ _1720_ _1721_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6140__B1 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_65_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8662__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ _1347_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8465__B _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _0316_ _0538_ _0620_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6097_ as2650.stack\[6\]\[12\] _1596_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5048_ _0334_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4284__I _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _1344_ _1304_ _2427_ _2428_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8738_ _0215_ clknet_leaf_41_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8669_ _0146_ clknet_leaf_7_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8499__A2 _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__A1 _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__A1 _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5843__I as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8120__A1 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8120__B2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4459__I _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5324__I3 as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6674__I _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5788__A3 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4922__I _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4748__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8535__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6849__I _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ _3928_ _3930_ _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8111__A1 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4281_ _3856_ _3861_ _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5476__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6020_ as2650.psl\[5\] _1535_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8716__D _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7971_ _2141_ _3936_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6976__A2 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6922_ _0429_ _2358_ _2353_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8178__A1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6853_ _2188_ _2256_ _2291_ _2295_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6728__A2 _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7925__A1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4832__I _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5804_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4739__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6784_ _2226_ _2227_ _1463_ _2173_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_52_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8523_ _0000_ clknet_leaf_76_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5735_ as2650.stack\[3\]\[7\] _1260_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8454_ _3767_ _3783_ _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5666_ _1138_ _1194_ _1218_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8350__A1 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5164__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7405_ _2817_ _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4617_ _4196_ _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8385_ as2650.psl\[5\] _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6900__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5597_ _4260_ _1156_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7336_ _2654_ _2753_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4548_ _3909_ _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8102__A1 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7267_ _2683_ net8 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_46_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _4059_ _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5467__A2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ _3985_ _1665_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7198_ _2595_ _2618_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8626__D _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ _1643_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8405__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6416__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6967__A2 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8169__A1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_55 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_66 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_77 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_88 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8558__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6719__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5838__I _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5942__A3 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__A1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4902__B2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6655__A1 _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5241__C _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7080__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A1 _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5630__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5394__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _1067_ _1103_ _1104_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8332__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7135__A2 _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_121_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5483__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6894__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4402_ as2650.ins_reg\[6\] _3983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8170_ _2844_ _0642_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5382_ _0519_ _0917_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7121_ as2650.stack\[7\]\[0\] _1019_ _2539_ _2542_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4333_ _3913_ _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7052_ _2434_ _3891_ _2468_ _2478_ _2479_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4264_ _3844_ _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _1511_ _1516_ _1519_ _1520_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__4827__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7203__I _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8399__A1 _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8700__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7071__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7954_ _1365_ _2603_ _2271_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_36_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6905_ _1348_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7885_ _3251_ _3264_ _3267_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6836_ _1054_ _1610_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6177__A3 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _0466_ _1975_ _2193_ _0727_ _2212_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_137_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ _2348_ _3829_ _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5718_ as2650.stack\[3\]\[0\] _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6698_ _1315_ _2152_ _1390_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8323__A1 _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7126__A2 _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8323__B2 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__B _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8437_ _1519_ _3766_ _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ as2650.stack\[0\]\[13\] _1066_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_80_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5688__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8368_ _3699_ _3703_ _3705_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7319_ _2734_ _2736_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7822__B _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8299_ _2997_ _3573_ _1708_ _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6637__A1 _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8209__I _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7113__I _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5860__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A1 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__B2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5568__I _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__B1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4472__I _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7365__A2 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8314__A1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5128__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8723__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5851__A2 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 io_in[7] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6862__I _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6800__A1 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4951_ _4209_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5478__I _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7670_ _3065_ _2582_ _3076_ _3077_ _2479_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4882_ _0466_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6621_ _1024_ _1045_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5367__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7693__I _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5906__A3 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6552_ _0796_ _2016_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8305__A1 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4965__I1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5503_ _1077_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6483_ _1952_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6867__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8222_ _0806_ _0802_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5434_ _1021_ _1012_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8153_ _3336_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5365_ _0941_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6619__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7104_ _2525_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4316_ _3895_ _3896_ _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8084_ _2333_ _3435_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5296_ _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7292__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6095__A2 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ _2461_ _2462_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5142__I1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8473__B _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6772__I _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7089__B _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7937_ as2650.stack\[7\]\[1\] _3294_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5388__I _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7868_ _1181_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6819_ _1057_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7799_ _3198_ _3199_ _3200_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6858__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8746__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5530__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7283__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__I _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5833__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7035__A1 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6682__I _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5597__A1 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5298__I _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7338__A2 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__I _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5150_ as2650.r0\[4\] _0366_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7274__A1 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6077__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ _0587_ _0605_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8724__D _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5588__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8771_ _0248_ clknet_leaf_55_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5983_ _1411_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7722_ _2276_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4934_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _0298_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7329__A2 _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7653_ _2727_ _2639_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4865_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6604_ _1004_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _2993_ _2994_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4796_ _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6535_ _1772_ _2011_ _2012_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8769__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4563__A2 _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _0611_ _1947_ _1658_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8468__B _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8205_ _2399_ _3548_ _3552_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5417_ _0845_ _0936_ _0933_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6397_ _1841_ _1842_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8136_ _3391_ _3485_ _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5348_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7265__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6068__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4287__I as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8067_ _0397_ _3349_ _3322_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5279_ as2650.psu\[2\] _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7018_ _3960_ _2073_ _2446_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5815__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7568__A2 _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5579__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8517__A1 _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7740__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7256__B2 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4490__A1 _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6767__B1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6231__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4650_ _3886_ _4229_ _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput10 wb_rst_i net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4581_ _4138_ _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6320_ _1713_ _1772_ _1773_ _1805_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6251_ _0784_ _1736_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5202_ _0699_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6182_ _4145_ _1659_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7247__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5133_ _0663_ _0669_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7798__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _0658_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4835__I _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A2 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8754_ _0231_ clknet_leaf_49_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5966_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6773__A3 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7705_ _4023_ _3111_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4917_ _0512_ _0514_ _0515_ _0418_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8685_ _0162_ clknet_leaf_7_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5981__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5897_ _1399_ _3963_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8591__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7636_ _0973_ _2875_ _3035_ _3045_ _3033_ _2620_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _0350_ _0442_ _0445_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6525__A3 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7567_ as2650.addr_buff\[2\] _2308_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4536__A2 _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _0295_ _0297_ _0300_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_88_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _0844_ _1758_ _1996_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7498_ _2863_ _2811_ _0712_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7486__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8629__D _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6449_ _1888_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8119_ _3463_ _3469_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5249__B1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7789__A2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6461__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6960__I _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__A2 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__A2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5972__A1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4480__I _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5724__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7477__A1 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__I _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7229__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7740__B _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4856__S _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5255__A3 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7966__I _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7401__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5820_ _1333_ _1334_ _1338_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5751_ _1237_ _1267_ _1274_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5963__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4702_ net7 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8470_ _3786_ _3798_ _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5682_ _1226_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7421_ _1639_ _2380_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4633_ _4212_ _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7352_ _2574_ _2767_ _2769_ _2739_ _2581_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4564_ _3874_ _4143_ _4144_ _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7468__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6303_ _1782_ _1787_ _1788_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7468__B2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7283_ as2650.addr_buff\[3\] _2152_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4495_ _3872_ _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6110__I _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6234_ _0767_ _0795_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6140__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6140__B2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6165_ _1651_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _1591_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8432__A3 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ _0555_ _0639_ _0640_ _0378_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_34_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8196__A2 _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8806_ _0283_ clknet_leaf_42_wb_clk_i as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7809__C _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6998_ _2355_ _1344_ _2387_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7943__A2 _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8737_ _0214_ clknet_leaf_43_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4757__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5949_ _1287_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8668_ _0145_ clknet_leaf_23_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__A2 _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5706__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7619_ as2650.pc\[12\] _0714_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8599_ _0076_ clknet_leaf_55_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5182__A2 _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7459__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8120__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6131__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4693__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7631__A1 _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4445__A1 _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7786__I _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8187__A2 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6198__A1 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__A2 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4748__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7698__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6122__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4280_ _3860_ _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6865__I _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7870__A1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7622__A1 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7970_ _2071_ _3324_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4436__A1 _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _1101_ _2356_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_54_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7696__I _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8178__A2 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _1503_ _2294_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7925__A2 _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5803_ _1029_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _1563_ _2078_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5936__A1 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4739__A2 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6105__I _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8522_ _3841_ _3842_ _1360_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5734_ _1244_ _1258_ _1262_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7689__A1 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8453_ _3769_ _3778_ _3781_ _3782_ _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5665_ as2650.stack\[1\]\[13\] _1135_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7404_ _2530_ _2818_ _2819_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8350__A2 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4616_ _4080_ _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5164__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8384_ _3671_ _1632_ _3716_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5596_ _1166_ _1074_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7335_ _1509_ _2600_ _2752_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4547_ net10 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8102__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7266_ _2683_ _2684_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4478_ _4057_ _4058_ _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6775__I _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6217_ _1657_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5467__A3 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7197_ _2587_ _2598_ _2610_ _2617_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6708__C _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ as2650.r123\[3\]\[0\] _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6416__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ _1127_ _1584_ _1588_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4427__A1 _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_56 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_67 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_78 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_89 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_109_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6015__I _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5942__A4 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6685__I as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7852__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7604__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7080__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__I _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5030__S _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7907__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6040__B1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6591__A1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8652__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8332__A2 _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5450_ _3959_ _1037_ _3880_ _3905_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_121_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6343__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4401_ _3913_ _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6894__A2 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5381_ _0937_ _0968_ _0970_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7120_ _2540_ _2541_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8096__A1 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4332_ as2650.ins_reg\[5\] _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8727__D _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7843__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7051_ _1358_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4263_ _3843_ _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4657__A1 _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6002_ _0396_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8399__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4409__A1 _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5004__I _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7953_ _2248_ _2261_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5939__I _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__I _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _2343_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7884_ as2650.stack\[4\]\[9\] _3266_ _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6835_ net25 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5909__A1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__A2 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6766_ as2650.r123\[2\]\[6\] _2197_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5717_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8505_ _3730_ _2347_ _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6697_ _1036_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8323__A2 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__C _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5648_ _1078_ _1189_ _1208_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6334__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8436_ _1451_ _2526_ _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8367_ net45 _3704_ _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6885__A2 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _0887_ _1010_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4896__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7318_ _2686_ _2735_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8298_ _2997_ _3617_ _2233_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6637__A2 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ as2650.stack\[5\]\[2\] as2650.stack\[4\]\[2\] _0883_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8525__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__A1 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__B2 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8011__A1 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6573__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5584__I _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8314__A2 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5128__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6876__A2 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8078__A1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4928__I _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5851__A3 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 io_in[8] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8250__A1 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _4074_ _0540_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6800__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8002__A1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4881_ _0467_ _0481_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6620_ _1026_ _1335_ _3904_ _1032_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_32_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6564__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__B2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5906__A4 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _1986_ _2002_ _2023_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5494__I _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8305__A2 _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5502_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6482_ _1953_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8221_ net51 _3567_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6867__A2 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5433_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8152_ _3408_ _3500_ _3501_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7642__C _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5364_ _0897_ as2650.stack\[1\]\[11\] as2650.stack\[0\]\[11\] _0901_ _0957_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_47_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8548__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7103_ _2180_ _1294_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4315_ as2650.cycle\[0\] _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6619__A2 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7816__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8083_ _2698_ _2177_ _3430_ _3434_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5295_ _0889_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7034_ _2109_ _2269_ _2236_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8698__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8241__A1 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4573__I _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7936_ _3285_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7867_ _3254_ _3249_ _3255_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6818_ _2240_ _2248_ _2261_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5358__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6555__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7817__C _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7752__B1 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7798_ _0528_ _3156_ _2790_ _0851_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6749_ _4127_ _2194_ _2198_ _2200_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6858__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8419_ _0362_ _0436_ _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__A1 _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5530__A2 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7807__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7124__I _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7283__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8480__A1 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7035__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8232__A1 _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5046__A1 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4483__I _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6794__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5597__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7743__B1 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8299__A1 _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__A4 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5080_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5489__I _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5037__A1 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6785__A1 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5588__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _1469_ _1476_ _1499_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8770_ _0247_ clknet_leaf_55_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4933_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7721_ _3101_ _3109_ _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4864_ _3957_ _0460_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7652_ _2105_ _3051_ _3059_ _3060_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_33_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6603_ _2064_ _2065_ _2067_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7583_ _1172_ _2967_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4795_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_59_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7209__I _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6113__I _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6534_ _0287_ _1656_ _2008_ as2650.r123_2\[1\]\[1\] _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5760__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6465_ _1940_ _1809_ _1945_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5952__I _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8204_ _2305_ _2399_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5416_ _1004_ _0967_ _0951_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7372__C _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6396_ _1794_ _1879_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5512__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8135_ _0616_ _0643_ _3484_ _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5347_ _0907_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7265__A2 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8066_ _0395_ _0390_ _3417_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5278_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8484__B _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7017_ _2306_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6776__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7919_ _3285_ _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6528__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8713__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5751__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6958__I _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8453__A1 _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8394__B _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6464__B1 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8205__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4490__A2 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6767__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6767__B2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4941__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7457__C _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7029__I _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7192__A1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _3992_ _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6250_ _0745_ _0790_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ _4108_ _0701_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6181_ _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8444__A1 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5132_ _0670_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5258__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _0659_ _0660_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_85_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4856__I1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5012__I _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7648__B _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6222__A3 _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8753_ _0230_ clknet_leaf_44_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5947__I _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5965_ _0711_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8736__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6773__A4 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7704_ _3110_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4916_ _4045_ _0412_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8684_ _0161_ clknet_3_3_0_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5896_ _1413_ _1059_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7635_ _2852_ _3036_ _3044_ _1636_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4847_ _0429_ _0447_ _0351_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7566_ _2974_ _2977_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4778_ _0377_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5733__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6930__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6517_ _0822_ _1759_ _1695_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7497_ _2823_ _2910_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _1928_ _1930_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5497__A1 _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4298__I _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6379_ _1520_ _1671_ _1862_ _1676_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8118_ _2916_ _1527_ _3467_ _3468_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_103_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7830__C _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8435__A1 _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8049_ _3332_ _3401_ _2647_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6997__A1 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6018__I _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6749__A1 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__A1 _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5972__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6921__A1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5724__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7477__A2 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5032__S0 _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8609__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7229__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7740__C _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8408__I _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5660__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8759__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__A2 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5750_ as2650.stack\[4\]\[3\] _1271_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5963__A2 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5681_ as2650.r123_2\[3\]\[6\] _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7165__A1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7420_ _2139_ _2604_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4632_ as2650.r0\[2\] _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6912__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8299__B _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7351_ _2768_ _2740_ _2470_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4563_ _3911_ _3947_ _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6302_ _0625_ _0471_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7468__A2 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7282_ _1347_ _2263_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4494_ _4065_ _4066_ _4071_ _4074_ _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6233_ _0767_ _0795_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6140__A2 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _3951_ _3850_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5115_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6095_ _1182_ _1592_ _1599_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5046_ _4122_ _0589_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8805_ _0282_ clknet_leaf_39_wb_clk_i as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6997_ _2426_ _2419_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5403__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_74_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5403__B2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4581__I _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8736_ _0213_ clknet_leaf_49_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _1458_ _1462_ _1465_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8667_ _0144_ clknet_leaf_24_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5879_ _1379_ _1382_ _1396_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7618_ _2975_ _3025_ _3027_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4509__A3 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5706__A2 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8598_ _0075_ clknet_leaf_31_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4530__B _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7549_ _0927_ _2875_ _2947_ _2960_ _2961_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8105__B1 _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6131__A2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__I0 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4756__I _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7631__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6971__I _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7735__C _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7698__A2 _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4381__A1 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4867__S _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6122__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7870__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7042__I _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7622__A2 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5633__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6881__I _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _2130_ _1532_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ _2083_ _1614_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7386__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5802_ _1312_ _1317_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_35_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6782_ _2225_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8521_ _2358_ _3833_ _3835_ _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7138__A1 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5733_ as2650.stack\[3\]\[6\] _1260_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6830__B _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7689__A2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8452_ _2160_ _1343_ _1329_ _1394_ _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5664_ _1138_ _1189_ _1217_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7403_ _0903_ as2650.stack\[3\]\[6\] as2650.stack\[2\]\[6\] _1014_ _1020_ _2819_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4615_ _4194_ _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5595_ _1165_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8383_ _3189_ _1630_ _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__I _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6900__A4 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7334_ _4144_ _2737_ _2739_ _2443_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4546_ _3993_ _4037_ _4126_ _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7265_ as2650.pc\[2\] as2650.pc\[1\] as2650.pc\[0\] _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4477_ _3909_ _3863_ _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5960__I _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7310__A1 _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6216_ _1679_ _1667_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7196_ _2612_ _2584_ _2613_ _2614_ _2616_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_131_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__A1 _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6147_ _1642_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ as2650.stack\[5\]\[6\] _1586_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4427__A2 _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6672__I0 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _0627_ _3860_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_57 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_68 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_79 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7377__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8719_ _0196_ clknet_leaf_38_wb_clk_i as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7127__I _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4363__A1 _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__I _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7852__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A2 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5863__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__I _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7604__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7368__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5918__A2 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__B2 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7540__A1 _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7037__I _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4400_ _3980_ _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5380_ _0882_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _3911_ _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8096__A2 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5780__I as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7050_ _2471_ _2477_ _2374_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4262_ as2650.ins_reg\[0\] _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_87_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7843__A2 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4657__A2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A1 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _1518_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4409__A2 _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7952_ net28 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6903_ _4009_ _2337_ _2342_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7359__A1 as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7883_ _1265_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6116__I _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6834_ net49 _2262_ _2275_ _2277_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5909__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6765_ _0649_ _2193_ _2210_ _2211_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5385__A3 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6582__A2 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5955__I _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4999__C _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8504_ _4225_ _3102_ _3818_ _3828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5716_ _1248_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4593__A1 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6696_ _2149_ _2150_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8435_ _3757_ _3764_ _3765_ _2435_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5647_ as2650.stack\[0\]\[12\] _1204_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6334__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__A1 _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8366_ _3681_ _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _0894_ _1012_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7317_ _2642_ _2643_ _2687_ _2690_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_85_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8087__A2 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4529_ _4109_ _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5690__I _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8297_ _2131_ _3620_ _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6098__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7248_ _0906_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7179_ _2599_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7598__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__A2 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8011__A2 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5865__I _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7770__A1 _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7522__A1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7522__B2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4336__A1 _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8078__A2 _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7825__A2 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__A2 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5836__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7589__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput9 io_in[9] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6261__A1 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4880_ _0478_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7210__B1 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5775__I _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__A2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6550_ as2650.r123_2\[1\]\[6\] _2015_ _2022_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5501_ _1082_ _1085_ _1087_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7990__I _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7513__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6481_ _1956_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8220_ _3566_ _3547_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5432_ _1019_ _0878_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8151_ net52 _3317_ _3472_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5363_ as2650.stack\[7\]\[11\] as2650.stack\[4\]\[11\] as2650.stack\[5\]\[11\] as2650.stack\[6\]\[11\]
+ _0884_ _0887_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__8069__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7102_ _1070_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4314_ as2650.cycle\[1\] _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8082_ _2214_ _2693_ _3431_ _3433_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5294_ _0877_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7033_ _2409_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__I _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6252__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7935_ _1228_ _3292_ _3297_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A2 _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7866_ as2650.stack\[5\]\[10\] _3252_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6004__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6817_ _2249_ _1618_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6555__A2 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7752__A1 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7797_ as2650.psl\[5\] _3113_ _0855_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5685__I _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7752__B2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4566__A1 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6748_ _2199_ _1756_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6679_ _3934_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8418_ _4194_ _3746_ _3748_ _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6858__A3 _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__A2 _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8349_ _1086_ _3685_ _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7807__A2 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5818__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4965__S _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8480__A2 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8642__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8232__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5046__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7440__B1 _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6794__A2 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7991__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5595__I _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6546__A2 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7743__A1 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__A1 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8299__A2 _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7743__C _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4939__I _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5809__A1 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8223__A2 _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5037__A2 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__C _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _1492_ _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6785__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7720_ _2448_ _4070_ _3125_ _3126_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_127_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4932_ as2650.r0\[5\] _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7651_ _2062_ _2630_ _3053_ _2635_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ _0462_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6537__A2 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7734__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ _0998_ _2032_ _2066_ _2054_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_127_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7582_ as2650.pc\[11\] _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4794_ _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _2001_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _3901_ _1691_ _1860_ _0643_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8203_ _2461_ _3533_ _3550_ _2316_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5415_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6395_ _0410_ _1837_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_28_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4720__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8134_ _3455_ _3482_ _3456_ _3483_ _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_5346_ as2650.stack\[7\]\[10\] as2650.stack\[4\]\[10\] as2650.stack\[5\]\[10\] as2650.stack\[6\]\[10\]
+ _0938_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7265__A3 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8065_ _3386_ _3415_ _3416_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ as2650.psu\[1\] _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7016_ _2300_ _2440_ _2444_ _2417_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8056__I _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__I _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6225__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6776__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7973__A1 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7918_ _3248_ _3284_ _3287_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4787__A1 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7849_ as2650.stack\[6\]\[4\] _3241_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4539__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8150__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A1 _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8453__A2 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8394__C _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A1 _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7661__B1 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__B2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8205__A2 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__A2 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7738__C _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__A2 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7192__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7754__B _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4950__A1 _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__I _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5200_ _4100_ _4104_ _4107_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_87_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6180_ _1666_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6884__I _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _0651_ _0672_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8444__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6455__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5258__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _4213_ _0469_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_opt_2_1_wb_clk_i_I clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7955__A1 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6758__A2 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8752_ _0229_ clknet_leaf_43_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _1296_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6222__A4 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7703_ _0443_ _0523_ _0863_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4915_ _0493_ _0386_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8683_ _0160_ clknet_leaf_17_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5895_ _1386_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6124__I _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7634_ _2885_ _3039_ _3043_ _2931_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4846_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8380__A1 _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ _2975_ _2976_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _4247_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_53_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6930__A2 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6516_ _0803_ _1860_ _1809_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7496_ as2650.pc\[7\] net2 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6447_ _1882_ _1886_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6143__B1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6694__A1 _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5497__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _0401_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8117_ _1108_ _3337_ _3126_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ _0904_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5249__A2 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6446__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8048_ _2893_ _3380_ _2650_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6997__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8199__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5421__A2 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5185__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6382__B1 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6921__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5032__S1 _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__A1 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5113__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A2 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5680_ _1225_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7165__A2 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7484__B _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4631_ _4210_ _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6912__A2 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__A1 _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7350_ _2572_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4562_ _4012_ _3944_ _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8114__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ as2650.r0\[7\] _0368_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7281_ _2698_ _2699_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4493_ _4073_ _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6676__A1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6232_ _1655_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6163_ _1650_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ as2650.stack\[6\]\[11\] _1596_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8703__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5100__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ _4201_ _0643_ _4118_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5651__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8050__B1 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8804_ _0281_ clknet_leaf_39_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6996_ _2391_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6282__C _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6600__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8735_ _0212_ clknet_leaf_55_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5947_ _1464_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8666_ _0143_ clknet_leaf_24_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5878_ _1383_ _1389_ _1391_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8353__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6789__I _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7617_ as2650.pc\[11\] _1488_ _3026_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4829_ _0429_ _0302_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_107_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8597_ _0074_ clknet_leaf_31_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5693__I _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_43_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4914__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7548_ _1366_ _2941_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8105__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7479_ _2396_ _2893_ _2851_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__I1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6029__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4525__S0 _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__I _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7147__A2 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8344__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4381__A2 _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5108__I _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5330__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__B2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6830__A1 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7479__B _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6383__B _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5778__I _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6850_ _2292_ _1311_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7386__A2 _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5801_ _1318_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5397__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6781_ _2075_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7993__I _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5936__A3 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8520_ _2357_ _3837_ as2650.psu\[3\] _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5732_ _1242_ _1258_ _1261_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8335__A1 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7138__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8451_ _2287_ _3779_ _3780_ _3781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5663_ as2650.stack\[1\]\[12\] _1213_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7689__A3 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7402_ _2624_ as2650.stack\[1\]\[6\] as2650.stack\[0\]\[6\] _2625_ _2818_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6897__A1 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4614_ _4169_ _4193_ _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8382_ _2916_ _1632_ _3715_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5594_ as2650.pc\[9\] _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_89_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7333_ as2650.addr_buff\[4\] _1416_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4545_ _4117_ _4125_ _3993_ _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5018__I _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7264_ as2650.pc\[3\] _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4476_ _3974_ _4056_ _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5462__B _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__I _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6215_ _3902_ _1664_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5321__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _2615_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6146_ _1384_ _1621_ _1630_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7074__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4507__S0 _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6077_ _1120_ _1584_ _1587_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6821__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6672__I1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input10_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_58 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_69 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7377__A2 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__C1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6979_ _2326_ _2224_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8718_ _0195_ clknet_leaf_36_wb_clk_i as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7836__C _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8326__A1 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8649_ _0126_ clknet_leaf_72_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8749__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4767__I _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7143__I _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7065__A1 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6812__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5615__A2 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__I _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4674__I0 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__C1 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5379__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5379__B2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__A2 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7746__C _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8317__A1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6879__A1 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5000__B1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7762__B _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7481__C _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4330_ as2650.ins_reg\[2\] _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4677__I _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ net26 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7053__I as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5854__A2 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7988__I _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7056__A1 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5067__B1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4409__A3 _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7951_ _1246_ _3286_ _3306_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _2341_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5301__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7882_ _3248_ _3264_ _3265_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7359__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4290__A1 _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6833_ _2276_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6031__A2 _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ as2650.r123\[2\]\[5\] _2197_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8308__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8503_ _3824_ _3827_ _1360_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5715_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5790__A1 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4593__A2 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _1038_ _1417_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8434_ _3727_ _3758_ _4023_ _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5646_ _1202_ _1182_ _1207_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4345__A2 _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8365_ _3700_ _1473_ _3702_ _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5971__I _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5577_ _1131_ _1144_ _1149_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8487__C _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7316_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4528_ _4108_ _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8296_ _3559_ _3639_ _3640_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7295__A1 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6098__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7247_ as2650.stack\[7\]\[2\] _0878_ _1019_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4459_ _4039_ _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7178_ _1051_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7047__A1 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6129_ _4139_ _1609_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6735__C _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7598__A2 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4536__B _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A2 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4281__A1 _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5211__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7770__A2 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8571__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5881__I _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__B _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7286__A1 _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7038__A1 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8235__B1 _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6217__I _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7249__S _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7210__A1 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6380__C _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7761__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5772__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5500_ _1086_ _1085_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6480_ _1959_ _1961_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5431_ _0876_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8150_ _1116_ _3409_ _3494_ _3499_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5362_ _0457_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7101_ _2522_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4313_ as2650.cycle\[5\] as2650.cycle\[4\] _3893_ _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8081_ _2175_ _2418_ _3432_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5293_ as2650.psu\[0\] _0886_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7032_ _3959_ _2438_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6252__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7934_ as2650.stack\[7\]\[0\] _3294_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7865_ _1174_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8594__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5966__I _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6004__A2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _2250_ _2251_ _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8342__I _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7796_ as2650.psu\[5\] _3138_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7752__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _4154_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5763__A1 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ _1535_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8498__B _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5629_ as2650.stack\[2\]\[13\] _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8417_ _4193_ _3747_ _4168_ _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__A3 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8348_ _3682_ _3687_ _3689_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7268__A1 as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8279_ _3602_ _3563_ _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5206__I _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__A2 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8480__A3 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6794__A3 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7991__A2 _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7577__B _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4780__I _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5754__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__A2 _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8201__B _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7259__A1 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5809__A2 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4955__I _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5980_ _1495_ _1496_ _0799_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4931_ _0523_ _0524_ _0528_ _0530_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7487__B _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5786__I _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4690__I as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7650_ _2768_ _3053_ _3058_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4862_ _3982_ _3887_ _4019_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6601_ _0997_ _2048_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7581_ _2966_ _2991_ _2992_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4793_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6532_ _1701_ _2002_ _2009_ _2010_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7498__A1 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _0986_ _1706_ _1944_ _1690_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8202_ _2327_ _3546_ _3549_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5414_ _0817_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6170__A1 _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6394_ _1876_ _1877_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8133_ _0542_ _0517_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5345_ _0886_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5026__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4720__A2 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8064_ _0305_ _0335_ _0336_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_102_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ as2650.psu\[0\] _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7015_ _2443_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_68_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4865__I _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7422__A1 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6225__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7917_ as2650.stack\[7\]\[8\] _3286_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4787__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7848_ _1103_ _3239_ _3243_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4539__A2 as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7779_ _3952_ _3114_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8150__A2 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A2 _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7661__A1 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7661__B2 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7151__I _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__A1 _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7754__C _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__A2 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8141__A2 _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5130_ _0652_ _0671_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7652__A1 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5061_ _0292_ _0367_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7996__I _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7404__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7955__A2 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4769__A2 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8751_ _0228_ clknet_leaf_44_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5963_ _1124_ _1479_ _1480_ _1450_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7010__B as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4914_ _0494_ _0513_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7702_ _3102_ _3107_ _3108_ _2299_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5894_ _1410_ _1411_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8682_ _0159_ clknet_leaf_73_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7633_ _2834_ _3030_ _3041_ _1607_ _3042_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _3981_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8380__A2 _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7664__C _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7564_ _2952_ _1157_ _0713_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ as2650.idx_ctrl\[1\] _3976_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_119_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6515_ _1003_ _1663_ _1994_ _1810_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7495_ _2777_ _2776_ _2908_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8132__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6446_ _0816_ _1186_ _1887_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6143__A1 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6143__B2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7680__B _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6694__A2 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8782__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6377_ _1669_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8116_ _2446_ _2737_ _3466_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5328_ _0920_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4595__I _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8047_ _3378_ _3380_ _3382_ _3319_ _3399_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6446__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5259_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4457__A1 _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7946__A2 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5957__A1 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__A3 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5709__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8371__A2 _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7574__C _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5185__A2 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6382__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7882__A1 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7634__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7634__B2 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__A1 _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7937__A2 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8655__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4620__A1 _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ _4073_ _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6373__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ _3902_ _3926_ _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8114__A2 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6300_ _1742_ _1749_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6125__A1 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7280_ _1068_ _3911_ _1092_ _1080_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_144_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7322__B1 _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4492_ _3988_ _4072_ _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6231_ as2650.r123_2\[2\]\[0\] _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6895__I _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6676__A2 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6162_ as2650.r123\[3\]\[7\] _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5113_ net2 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7625__A1 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _1175_ _1592_ _1598_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5487__I0 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5100__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__B _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6336__S _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7928__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8050__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8803_ _0280_ clknet_3_1_0_wb_clk_i as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8050__B2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _2417_ _2420_ _2423_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6135__I _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8734_ _0211_ clknet_leaf_55_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5946_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4611__A1 _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8665_ _0142_ clknet_leaf_23_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5877_ _1392_ _4072_ _1394_ _4207_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7616_ _3005_ _2976_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4828_ as2650.holding_reg\[3\] _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8596_ _0073_ clknet_leaf_54_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7547_ _2951_ _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4759_ _0356_ _0360_ _3998_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8105__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7478_ _2599_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7864__A1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6429_ _1655_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4678__A1 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_12_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8528__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7616__A1 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__S1 _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8678__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4850__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6355__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4721__C _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6107__A1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7855__A1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4669__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8280__A1 _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8032__A1 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ _3920_ _3995_ _3932_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_35_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6780_ _2108_ _3929_ _2073_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_35_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6594__A1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5397__A2 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5731_ as2650.stack\[3\]\[5\] _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5794__I _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8335__A2 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8450_ _4135_ _1410_ _2675_ _2335_ _2512_ _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5149__A2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5662_ _1211_ _1182_ _1216_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7689__A4 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7401_ _2530_ _2815_ _2816_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4613_ _4173_ _4192_ _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6897__A2 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8381_ _2130_ _1630_ _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5593_ _1155_ _1162_ _1164_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7332_ _2746_ _2748_ _2749_ _2661_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4544_ _4119_ _4124_ _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6649__A2 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7846__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7263_ _2581_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _3888_ _3984_ _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5857__B1 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6214_ _1656_ _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5462__C _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7194_ _1615_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5321__A2 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _1563_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7074__A2 _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8271__A1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ as2650.stack\[5\]\[5\] _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4507__S1 _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6821__A2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _0625_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8023__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_59 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6034__B1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6034__C2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6978_ _2374_ _1313_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8717_ _0194_ clknet_leaf_33_wb_clk_i as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8648_ _0125_ clknet_leaf_71_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7534__B1 _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5209__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8579_ _0056_ clknet_leaf_61_wb_clk_i as2650.r123_2\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7837__A1 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7065__A2 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8262__A1 _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4823__A1 _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4674__I1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8014__A1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6025__B1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__C2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8317__A2 _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6328__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__B2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6879__A2 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5000__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5551__A2 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7828__A1 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6500__A1 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A3 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8253__A1 _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8253__B2 _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__I _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5067__A1 _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__B2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7950_ as2650.stack\[7\]\[7\] _3283_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4814__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8005__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6901_ _1379_ _1382_ _2254_ _4056_ _2340_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7881_ as2650.stack\[4\]\[8\] _1277_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4290__A2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6832_ _1357_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _4155_ _1965_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8502_ _2358_ _3826_ _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6319__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5714_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6694_ _3941_ _2147_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5790__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8433_ _3763_ _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5645_ as2650.stack\[0\]\[11\] _1204_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4345__A3 _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5576_ as2650.stack\[1\]\[7\] _1146_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8364_ _1109_ _3701_ _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5473__B _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7315_ as2650.pc\[4\] net9 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4868__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4527_ _4100_ _4104_ _4107_ _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7819__A1 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8295_ net38 _3557_ _3614_ _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8492__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4458_ _4038_ _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7246_ _2549_ _2649_ _2665_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7177_ _2596_ _2597_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4389_ _3969_ _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7047__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6128_ _1516_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6059_ _1574_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4281__A2 _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6558__A1 _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8716__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5781__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6730__A1 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8483__A1 _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8235__A1 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7038__A2 _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8235__B2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6797__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6549__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7757__C _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7210__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5221__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5772__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ as2650.psu\[2\] _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ as2650.r123\[0\]\[3\] _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4312_ _3891_ _3892_ _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7100_ _2272_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8080_ _2881_ _3414_ _2703_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8474__A1 _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5292_ as2650.stack\[7\]\[8\] as2650.stack\[4\]\[8\] as2650.stack\[5\]\[8\] as2650.stack\[6\]\[8\]
+ _0885_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7031_ _2434_ _1037_ _2435_ _2459_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6788__A1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5312__I _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4638__I1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7933_ _3262_ _3292_ _3296_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8739__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7864_ _3251_ _3249_ _3253_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _0458_ _0853_ _2257_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__5212__A1 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7795_ _3143_ _0805_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5212__B2 _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ as2650.r123\[2\]\[0\] _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5763__A2 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6677_ _2133_ _2120_ _2135_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8416_ _3745_ _4036_ _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5628_ _1154_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5915__C _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8347_ net41 _3688_ _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5559_ as2650.stack\[1\]\[0\] _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7268__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8278_ _1166_ _1159_ _1485_ _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5931__B _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _1092_ _2589_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7976__B1 _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7440__A2 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6794__A4 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6951__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5754__A2 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__A3 _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6988__I _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5892__I _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6703__A1 _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6937__B _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5809__A3 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8208__A1 _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8208__B2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7431__A2 _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4930_ _0529_ _0521_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _3967_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6600_ _1985_ _2027_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4792_ net8 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7580_ _2276_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6942__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6531_ _4153_ _4158_ _1912_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4953__B1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7498__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6462_ _0614_ _1680_ _1943_ _1706_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8111__C _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8201_ _3366_ _3548_ _2465_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5413_ as2650.r123\[0\]\[7\] _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6393_ _1836_ _1844_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6170__A2 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8447__A1 _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5344_ _0885_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8132_ _0541_ _0517_ _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6847__B _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5275_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8063_ _0335_ _0336_ _0306_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_138_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7014_ _2442_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8561__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__I _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7678__B _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5977__I _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7916_ _3285_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_37_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__A3 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4814__C _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7186__A1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7847_ as2650.stack\[6\]\[3\] _3241_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5736__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7778_ _3178_ _3179_ _2316_ _3180_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5292__S0 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _2180_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4711__A3 _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7110__B2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7661__A2 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__A2 _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7588__B _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4791__I _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7770__C _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8429__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8584__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4966__I _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5060_ _4079_ _0566_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7404__A2 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__I _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8750_ _0227_ clknet_leaf_52_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _1479_ _1461_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7701_ _2344_ _4203_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4913_ _0310_ _0328_ _0381_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8681_ _0158_ clknet_leaf_73_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5893_ _3946_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7632_ _2611_ _3033_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ _0444_ _0303_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5718__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7563_ _2944_ _2942_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_53_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4775_ _4160_ _0364_ _0376_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7517__I _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6514_ _0804_ _1683_ _1992_ _1993_ _1662_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7494_ _2825_ _2829_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6445_ _1926_ _1927_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6143__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6376_ _1686_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7891__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8115_ _3332_ _3465_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5327_ _0921_ as2650.stack\[1\]\[9\] as2650.stack\[0\]\[9\] _0901_ _0922_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_142_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8046_ _3321_ _3398_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ _0851_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4457__A2 _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5189_ _4212_ _0526_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8199__A3 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5406__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A2 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7159__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5709__A2 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6906__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4917__B1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6382__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7331__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7882__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__C _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7634__A2 _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7398__A1 _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8207__B _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5948__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4620__A2 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7765__C _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7570__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4560_ _4140_ _3931_ _3937_ _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_50_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4384__A1 as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4491_ _3940_ _3919_ _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7322__A1 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6125__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7322__B2 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6230_ _1716_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7873__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5884__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4696__I _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6161_ _1649_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _0627_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ as2650.stack\[6\]\[10\] _1596_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5636__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__I1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _0512_ _0639_ _0640_ _0418_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7389__A1 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8117__B _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__B _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8802_ _0279_ clknet_leaf_41_wb_clk_i as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8050__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _1312_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8733_ _0210_ clknet_leaf_54_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _1376_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8664_ _0141_ clknet_leaf_21_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5876_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7615_ _2973_ _3004_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4827_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7561__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8595_ _0072_ clknet_leaf_32_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4375__A1 _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7546_ _2588_ _2953_ _2954_ _2958_ _2446_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4758_ _0357_ _0340_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7313__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7477_ _2437_ _2890_ _2891_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5990__I _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4689_ _4185_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6428_ as2650.r123_2\[2\]\[4\] _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7864__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5875__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__A2 _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6359_ _1839_ _1843_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7616__A2 _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8029_ _2644_ _3381_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_52_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7092__A3 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4850__A2 _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6052__A1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8329__B1 _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A2 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7157__I _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7552__A1 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4366__A1 as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6996__I _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7304__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7855__A2 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A2 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__A2 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8622__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8032__A2 _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6043__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7776__B _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7791__A1 _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8772__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5730_ _1251_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8335__A3 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ as2650.stack\[1\]\[11\] _1213_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7543__A1 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7400_ as2650.stack\[6\]\[6\] _1014_ _0890_ as2650.stack\[7\]\[6\] _0879_ _2816_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4612_ _4179_ _4188_ _4191_ _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8380_ _3699_ _3713_ _3714_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5592_ as2650.stack\[2\]\[8\] _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7331_ _1508_ _2551_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4543_ _4123_ _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4420__S _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7846__A2 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7262_ _2521_ _2680_ _2681_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4474_ _4054_ _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7016__B _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5857__B2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _4037_ _1658_ _1694_ _1699_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7193_ _1030_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5321__A3 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _1640_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8271__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _1577_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__A1 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5026_ as2650.r0\[6\] _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6034__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6034__B2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _2373_ _2407_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5985__I _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__B _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7782__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8361__I _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4596__A1 _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8716_ _0193_ clknet_leaf_32_wb_clk_i as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5928_ _0826_ _0837_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5918__C _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8647_ _0124_ clknet_3_1_0_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5859_ _1308_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6337__A2 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7534__B2 _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8578_ _0055_ clknet_leaf_62_wb_clk_i as2650.r123_2\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5934__B _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7529_ _1165_ _0712_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7298__B1 as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7837__A2 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5848__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5225__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8645__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8262__A2 _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8795__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8014__A2 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6025__B2 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5895__I _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7773__A1 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6328__A2 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6005__B _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7525__A1 _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6879__A3 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5000__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7828__A2 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6500__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7350__I _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4814__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _3986_ _2252_ _2338_ _2339_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_76_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8005__A2 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7880_ _1268_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6016__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6831_ _2268_ _2274_ _2262_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__A1 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6762_ _0560_ _2193_ _2208_ _2209_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8501_ _3730_ _3825_ _3819_ _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5713_ _1133_ _1152_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6693_ _1389_ _1391_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7516__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6319__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8432_ _3727_ _3758_ _3762_ _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5644_ _1202_ _1175_ _1206_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8363_ _3683_ _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8130__B _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5575_ _1127_ _1144_ _1148_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7314_ _2731_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4526_ _4105_ _4106_ _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4750__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7819__A2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8294_ _2965_ _3409_ _3638_ _3374_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7245_ _2418_ _2655_ _2664_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8492__A2 _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4457_ _3987_ _3938_ _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4502__A1 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _1080_ _1514_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4388_ as2650.ins_reg\[2\] as2650.ins_reg\[3\] _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _0849_ _1621_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8244__A2 _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6058_ _1011_ _1017_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _0433_ _0594_ _0598_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8305__B _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6558__A2 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__A1 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__A1 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6604__I _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5230__A2 _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7507__A1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8180__A1 _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8483__A2 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4794__I _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8235__A2 _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6797__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6549__A2 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5221__A2 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5360_ _0932_ _0934_ _0953_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4311_ as2650.cycle\[2\] _3892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5291_ _0886_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__A1 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7030_ _2449_ _2455_ _2457_ _2458_ _2164_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8226__A2 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7985__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6788__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7985__B2 _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__A1 _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7932_ as2650.stack\[7\]\[14\] _3294_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7863_ as2650.stack\[5\]\[9\] _3252_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _3879_ _1054_ _1615_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_51_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7794_ _1464_ _0622_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5212__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6745_ _2196_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4971__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ _2134_ _2126_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8162__A1 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8415_ _3745_ _4036_ _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5627_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8346_ _3681_ _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4723__A1 _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _4083_ _4086_ _4089_ _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8277_ _2128_ _3619_ _3621_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5489_ _1065_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6476__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7228_ _2639_ _2638_ _2647_ _2346_ _2392_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7159_ _2521_ _2577_ _2580_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6228__A1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__A2 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7976__A1 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7976__B2 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8035__B _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5203__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6951__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4789__I _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6703__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_7_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5841__C _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8208__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5413__I as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4860_ _3972_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8392__A1 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _0312_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6942__A2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6530_ as2650.r123_2\[1\]\[0\] _2008_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4953__A1 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8144__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6461_ _0804_ _1668_ _1942_ _1761_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7075__I _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8200_ net35 _3547_ _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5412_ _0990_ _0934_ _1001_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6392_ _1839_ _1843_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8131_ _3350_ _3479_ _3480_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5343_ _0910_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_142_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8447__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8062_ net31 _3413_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5274_ _0851_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7024__B _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7013_ _2421_ _1399_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8706__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__I _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7958__A1 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6630__A1 _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7915_ _3282_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7846_ _1097_ _3239_ _3242_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7186__A2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8383__A1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_77_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7777_ _3164_ _0511_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5993__I _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4989_ _0531_ _0535_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6728_ _1384_ _3945_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5292__S1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4944__A1 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8135__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6146__B1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6659_ _2121_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4402__I as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8329_ _3661_ _3666_ _3670_ _3671_ _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_106_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8438__A2 _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7713__I _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4711__A4 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7949__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6621__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8374__A1 _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__B2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5408__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6688__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8429__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5143__I _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6860__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5663__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5961_ _1284_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_3_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7700_ _3050_ _4037_ _3106_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4912_ _0417_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8680_ _0157_ clknet_leaf_2_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__S _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5892_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8365__A1 _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7168__A2 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7631_ _2749_ _3040_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4843_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8403__B _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__S _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7562_ _2973_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8117__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ as2650.r123\[1\]\[2\] _4253_ _0375_ _4154_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ _0813_ _1682_ _1703_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7493_ as2650.pc\[8\] _0711_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _1920_ _1925_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5351__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _1807_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8114_ _2133_ _2881_ _3464_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5326_ _0896_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8045_ _3348_ _3390_ _3397_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5257_ _4184_ _0463_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_69_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7643__A3 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6851__A1 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5188_ _4079_ _0744_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5988__I _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5957__A3 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5002__B _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7829_ as2650.psu\[7\] _3114_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6906__A2 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4917__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4917__B2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5228__I _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7331__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7095__A1 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6842__A1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5645__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8207__C _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6008__B _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6070__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4307__I _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8347__A1 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A1 _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7570__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4384__A2 as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7781__C _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ _3950_ _4070_ _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__A2 _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6125__A3 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5884__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6160_ as2650.r123\[3\]\[6\] _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7086__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5111_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6091_ _1169_ _1592_ _1597_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5636__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5042_ _4045_ _0589_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7389__A2 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8801_ _0278_ clknet_leaf_65_wb_clk_i as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6993_ _2421_ _2281_ _2411_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8732_ _0209_ clknet_leaf_54_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5944_ _1420_ _1461_ _1349_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8663_ _0140_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5875_ _1043_ _3910_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4661__B _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7010__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4826_ as2650.holding_reg\[3\] _0302_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7614_ _1185_ _2772_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8594_ _0071_ clknet_leaf_32_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7561__A2 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4375__A2 _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7545_ _2444_ _2941_ _2957_ _1317_ _2701_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4757_ _0358_ _0341_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7476_ _2888_ _2847_ _2889_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4688_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7313__A2 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8510__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6427_ _1716_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6521__B1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7263__I _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5875__A2 _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__A3 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6358_ _1841_ _1842_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5309_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6289_ _1722_ _1755_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6824__A1 _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8028_ _3345_ _2640_ _2641_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5511__I _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_21_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8329__B2 _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7438__I _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7001__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7882__B _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8501__A1 _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5315__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__I _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_opt_2_0_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4669__A3 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8265__B1 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6815__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8017__B1 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6291__A2 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__A2 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7791__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _1211_ _1175_ _1215_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7543__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _4028_ _4190_ _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4357__A2 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5554__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5591_ _1154_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7330_ _2377_ _2747_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4542_ _4032_ _4122_ _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5306__A1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7261_ _1093_ _2578_ _2579_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4473_ _4053_ _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5306__B2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5857__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4500__I _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6212_ _1695_ _1698_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7016__C _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7192_ _2215_ _2598_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7059__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _1325_ _1621_ _1632_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7811__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6806__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6074_ _1112_ _1584_ _1585_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5025_ _0618_ _4228_ _0623_ _4211_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8597__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7231__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6034__A2 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6976_ _2374_ _2375_ _1338_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7782__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8715_ _0192_ clknet_leaf_33_wb_clk_i as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5927_ _1443_ _0830_ _1444_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6990__B1 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5858_ _1048_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8646_ _0123_ clknet_leaf_73_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7534__A2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ _1007_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8577_ _0054_ clknet_3_4_0_wb_clk_i as2650.r123_2\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7528_ _1165_ _2940_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7298__A1 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7298__B2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7459_ _0881_ _2870_ _2873_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5506__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4566__B _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__A2 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__I _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7525__A2 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6879__A4 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8501__B _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7289__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__I0 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7461__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5472__B1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6016__A2 _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7213__A1 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6830_ _2096_ _2270_ _2273_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5224__B1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6761_ as2650.r123\[2\]\[4\] _2202_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4578__A2 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6972__B1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8500_ _0962_ _2356_ _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5712_ _1246_ _1240_ _1247_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5643_ as2650.stack\[0\]\[10\] _1204_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8431_ _3153_ _4203_ _3761_ _1504_ _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8411__B _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5527__S _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6710__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8362_ _3683_ _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5574_ as2650.stack\[1\]\[6\] _1146_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7313_ _1347_ _2249_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4525_ as2650.r123\[1\]\[7\] as2650.r123\[0\]\[7\] as2650.r123_2\[1\]\[7\] as2650.r123_2\[0\]\[7\]
+ _3845_ _3856_ _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8293_ _3622_ _3632_ _3637_ _1465_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4750__A2 _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5326__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7244_ _2659_ _2660_ _2662_ _2663_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _4036_ _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8492__A3 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7175_ as2650.pc\[0\] net5 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4502__A2 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4387_ _3967_ _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ _1621_ _1623_ _1624_ _1626_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7452__A1 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6057_ _1264_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5008_ _4015_ _0600_ _0602_ _0350_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5996__I _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6558__A3 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__A2 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A2 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5766__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _2385_ _1390_ _2388_ _2389_ _2375_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_74_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4405__I _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8629_ _0106_ clknet_leaf_12_wb_clk_i as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7716__I _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8180__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6191__A1 _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7691__A1 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8762__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7746__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4315__I as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8171__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6182__A1 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5146__I _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4310_ as2650.cycle\[3\] _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7131__B1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5290_ as2650.psu\[1\] _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7682__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6485__A2 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4496__A1 _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7985__A2 _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4638__I3 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7931_ _3260_ _3292_ _3295_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__A2 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6705__I _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7310__B _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7862_ _1574_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6813_ _2256_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7793_ _3164_ _0611_ _3168_ _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5212__A3 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6744_ _4128_ _4136_ _2195_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_56_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ as2650.addr_buff\[4\] _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4971__A2 _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8162__A2 _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5626_ _1191_ _1179_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8414_ _4027_ _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6173__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8785__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5557_ _1134_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5920__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8345_ _3684_ _4203_ _3686_ _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4723__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4508_ _4087_ _4088_ _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_8276_ _3591_ _3620_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6476__A2 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7227_ _2422_ _2646_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4439_ _4019_ _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ _2524_ _2578_ _2579_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6109_ _1052_ _1045_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7425__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__A2 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7089_ _1035_ _2081_ _2103_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7976__A2 _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5987__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7728__A2 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6400__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4411__A1 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6164__A1 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7900__A2 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__A1 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__A1 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6467__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4478__A1 _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7416__A1 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5978__A1 _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8658__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8392__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4790_ _0294_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4953__A2 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8144__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6460_ _0622_ _1812_ _1941_ _1762_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5411_ _0991_ _0858_ _0869_ _1000_ _0861_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6391_ _1873_ _1874_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5902__A1 _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8130_ _0618_ _3354_ _3348_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5342_ _0858_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8061_ net30 net29 net28 _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7655__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5273_ _0868_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7091__I _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4469__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7012_ _2142_ _2436_ _2281_ _2440_ _2264_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7024__C _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7407__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7958__A2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8080__A1 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6630__A2 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7914_ _3283_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7845_ as2650.stack\[6\]\[2\] _3241_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8383__A2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7776_ _2492_ _0557_ _3050_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4988_ _0586_ _0538_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6727_ _2179_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4944__A2 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8135__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6146__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ as2650.addr_buff\[0\] _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6146__B2 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5609_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ as2650.r123_2\[0\]\[4\] _2044_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_139_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8328_ _3080_ _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__B _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7646__A1 as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8259_ _2410_ _3604_ _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5514__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5121__A2 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7949__A2 _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8071__A1 _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6621__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8374__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A2 _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8126__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6137__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7334__B1 _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6688__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7885__A1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7637__A1 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__I _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6860__A2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8062__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ _1477_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5891_ _3875_ _3910_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8365__A2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7630_ as2650.addr_buff\[4\] _2384_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4842_ _3972_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8403__C _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7561_ as2650.pc\[10\] _1487_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4773_ _4258_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8117__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6512_ _0807_ _1671_ _1991_ _1676_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7492_ _2781_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _1920_ _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6374_ _1806_ _1822_ _1823_ _1858_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8113_ _2377_ _3446_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5325_ _0907_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5103__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ _3846_ _0522_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8044_ _1518_ _3391_ _3396_ _2401_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__A2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5187_ _0774_ _0782_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__A1 _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8053__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5957__A4 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8356__A2 _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7828_ _0810_ _1625_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7759_ _1094_ _3100_ _3163_ _3129_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8108__A2 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6119__A1 _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7867__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7724__I _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7619__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7095__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8292__A1 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8292__B2 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6784__B _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8044__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6075__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8504__B _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5419__I _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4323__I _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4384__A3 as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _0419_ _0682_ _0703_ _0512_ _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__7086__A2 _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ as2650.stack\[6\]\[9\] _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5097__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _0537_ _0620_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4844__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8035__A1 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8800_ _0277_ clknet_leaf_9_wb_clk_i as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6597__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6992_ _1614_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6597__B2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8731_ _0208_ clknet_leaf_53_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5943_ _1459_ _1460_ _0817_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8338__A2 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6713__I _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8662_ _0139_ clknet_leaf_69_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5874_ _1308_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__C _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7010__A2 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _3022_ _3023_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4825_ _4165_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8593_ _0070_ clknet_leaf_34_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5329__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7544_ _2605_ _2956_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5572__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ _4028_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7475_ _2888_ _2847_ _2889_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4687_ _4214_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8510__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6426_ _1859_ _1908_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__A1 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__B2 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4532__B1 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6357_ _0533_ _0527_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7077__A2 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6288_ _1725_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5088__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5999__I _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8027_ net30 _3379_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6824__A2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _0824_ _0596_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8026__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5948__B _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7719__I _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8719__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7001__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_72_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_61_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4366__A3 _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6760__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6498__C _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6512__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8265__A1 _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6815__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8017__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4429__I1 _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5003__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _4163_ _4189_ _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7792__C _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5590_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4357__A3 _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5554__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ _4120_ _4121_ _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4762__B1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7364__I _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4472_ _4000_ _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6503__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7260_ _2523_ _2677_ _2679_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6201__C _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6211_ _4124_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7191_ _2611_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6142_ _1550_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6806__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ as2650.stack\[5\]\[4\] _1580_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4429__S _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__C _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8008__A1 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _4228_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7231__A2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ _1465_ _2395_ _2404_ _2405_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5242__A1 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8714_ _0191_ clknet_leaf_30_wb_clk_i as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5926_ _0695_ _0685_ _0829_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6990__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6990__B2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8645_ _0122_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5857_ _1363_ _1367_ _1370_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8576_ _0053_ clknet_leaf_67_wb_clk_i as2650.r123_2\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5788_ _4135_ _0855_ _1058_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6599__B _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ _2937_ _2902_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4739_ _0339_ _4221_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_120_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8495__A1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7458_ _2757_ _2871_ _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7207__C _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ _1829_ _1891_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7389_ _2675_ _2790_ _2805_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__B _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5522__I as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8541__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7449__I _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6733__A1 _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7289__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8238__A1 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8229__B _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7461__A2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5472__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5472__B2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__A3 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8410__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7213__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5224__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5224__B2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6760_ _4155_ _1938_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6972__A1 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4578__A3 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6972__B2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5711_ as2650.stack\[2\]\[7\] _1229_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6691_ _4129_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8430_ _1531_ _1457_ _3760_ _3153_ _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5642_ _1202_ _1169_ _1205_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8361_ _3681_ _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5573_ _1120_ _1144_ _1147_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4511__I _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7312_ _1106_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4524_ _4087_ _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8477__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8292_ _2965_ _3495_ _3636_ _2595_ _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7243_ _1517_ _2603_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4455_ _3998_ _4011_ _4031_ _4035_ _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_67_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7174_ _2303_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4386_ _3861_ _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8564__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6125_ _1625_ _1337_ _1620_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5342__I _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _1426_ _1571_ _1572_ _1359_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5007_ _0603_ _0605_ _0354_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8401__A1 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5215__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _1383_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6963__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5766__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _1361_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6889_ _2144_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8628_ _0105_ clknet_3_2_0_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6715__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8559_ _0036_ clknet_leaf_43_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6191__A2 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4421__I _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8468__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7140__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7732__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7140__B2 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8049__B _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5252__I _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7443__A2 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5454__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7400__C _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7179__I _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5757__A2 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5509__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6182__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4331__I _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8459__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6967__B _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8587__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7131__A1 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7131__B2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7682__A2 _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4496__A2 _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7930_ as2650.stack\[7\]\[13\] _3294_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ _1168_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7198__A1 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ _2252_ _2254_ _2255_ _1406_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_58_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6922__S _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6945__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5748__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7792_ _2323_ _1940_ _3193_ _2399_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6743_ _2192_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4956__B1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4956__C2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6721__I _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6674_ _1541_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7038__B _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8413_ _0362_ _0436_ _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5625_ _0528_ _1073_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7370__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6173__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4803__S0 _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7370__B2 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8344_ _1072_ _3685_ _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5556_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4507_ as2650.r123\[1\]\[1\] as2650.r123\[0\]\[1\] as2650.r123_2\[1\]\[1\] as2650.r123_2\[0\]\[1\]
+ _3857_ _3854_ _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_69_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8275_ _2997_ _3617_ _3618_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5487_ _1071_ _1072_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7226_ _2421_ _2645_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _3983_ _3916_ _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7157_ _2167_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4369_ _3949_ _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6108_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7088_ _2507_ _2508_ _2509_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _1514_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5987__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__A1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7727__I _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4411__A2 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7361__A1 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__A2 _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6703__A4 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4478__A2 _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5427__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8507__B _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5710__I _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5978__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4650__A2 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8392__A3 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7352__A1 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7352__B2 _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _0867_ _0997_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6390_ _1853_ _1856_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5902__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5341_ _0364_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8060_ _2688_ _3411_ _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7655__A2 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5272_ _4131_ _0856_ _0465_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4469__A2 _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5666__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7011_ _2437_ _2438_ _2439_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_114_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7407__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8417__B _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6466__I0 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7958__A3 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8080__A2 _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6091__A1 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8602__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout51_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7913_ _3282_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6630__A3 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7844_ _1590_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7775_ _2486_ _0518_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8752__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ as2650.holding_reg\[5\] _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6726_ _4076_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6657_ _2119_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6146__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5608_ as2650.pc\[11\] _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7894__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6588_ _2052_ _2055_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8327_ _1185_ _3502_ _3669_ _3031_ _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5539_ as2650.stack\[0\]\[5\] _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4839__C _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8258_ _2943_ _3563_ _3602_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7646__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _2528_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_15_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8189_ _3383_ _3536_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5409__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6626__I _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6082__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__A1 _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6137__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7334__B2 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7885__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5896__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7637__A2 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4320__A1 _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8625__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8775__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5820__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4910_ _0490_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5890_ _1371_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _0432_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7573__A1 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _1172_ _2971_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4772_ _0370_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_92_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6511_ _0810_ _1861_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7325__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7491_ _2775_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6442_ _1923_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7876__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5887__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6373_ _1719_ _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8112_ _3132_ _3462_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5324_ as2650.stack\[7\]\[9\] as2650.stack\[4\]\[9\] as2650.stack\[5\]\[9\] as2650.stack\[6\]\[9\]
+ _0885_ _0887_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7628__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5639__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8043_ _3391_ _3395_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5255_ _3994_ _0462_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5103__A3 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5186_ _0408_ _0562_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4862__A2 _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6890__B _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5811__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7827_ _3131_ _0844_ _3225_ _3226_ _3149_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7564__A1 _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7277__I _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6181__I _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7758_ _3152_ _3161_ _3162_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6709_ _3953_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7689_ _2092_ _2218_ _3094_ _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_123_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7867__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5878__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4925__I0 as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5525__I _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8648__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4550__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7619__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8292__A2 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6784__C _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4302__A1 _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8798__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4853__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8044__A2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5260__I _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__S _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__I _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7915__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6959__C _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5869__A1 _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6530__A2 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7086__A3 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5097__A2 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _0537_ _0619_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4844__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6991_ _1024_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6597__A2 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7794__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8730_ _0207_ clknet_leaf_51_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5942_ _0710_ _0613_ _0410_ _0391_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_80_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8661_ _0138_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5873_ _3903_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7546__A1 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7546__B2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4514__I _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7612_ _1178_ _2809_ _2191_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4824_ _4119_ _0390_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8592_ _0069_ clknet_leaf_34_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5021__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7543_ _2955_ _2309_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4755_ _4021_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7474_ net3 _4103_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7849__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4686_ _4160_ _4252_ _0288_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6425_ _1758_ _1906_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8510__A3 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6521__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6356_ _1838_ _1840_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4532__B2 _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5307_ _0875_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8274__A2 _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6287_ as2650.r123_2\[2\]\[1\] _1717_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6285__A1 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5088__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8026_ net53 net28 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _0828_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8026__A2 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5169_ _0738_ _0758_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5080__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6588__A2 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7785__A1 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__A1 _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7537__A1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6760__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_30_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6512__A2 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4523__A1 _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8265__A2 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7470__I _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5079__A2 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7403__C _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6086__I _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4826__A2 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8017__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__A2 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7776__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7528__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4334__I as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ as2650.idx_ctrl\[1\] _3976_ _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4762__B2 _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ _4051_ _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6503__A2 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7700__A1 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6210_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7190_ _1633_ _1322_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _1626_ _1637_ _1638_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6806__A3 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _1575_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5023_ _0593_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6019__A1 _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7767__A1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8425__B _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6724__I _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6974_ _1527_ _1327_ _2184_ _1504_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5925_ as2650.psl\[1\] _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8713_ _0190_ clknet_leaf_30_wb_clk_i as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7519__A1 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6990__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8644_ _0121_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ _0464_ _4164_ _1371_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8192__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4807_ as2650.r0\[4\] _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8798__D _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8575_ _0052_ clknet_leaf_46_wb_clk_i as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5787_ _0840_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4753__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7526_ _2521_ _2936_ _2939_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4738_ _0339_ _4221_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7457_ _0904_ as2650.stack\[3\]\[7\] as2650.stack\[2\]\[7\] _2668_ _1021_ _2872_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4669_ _4202_ _4092_ _4248_ _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8495__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _1831_ _1845_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7388_ _2635_ _2774_ _2804_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7504__B _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6339_ _1786_ _1799_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5803__I _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8009_ net53 _3307_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4419__I _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7758__A1 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6634__I _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8054__C _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6981__A2 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8183__A1 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6733__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6497__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5544__I0 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8238__A2 _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6249__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7997__A1 _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4329__I _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5472__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8410__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6421__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6972__A2 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5710_ _1130_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6690_ _1423_ _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8174__A1 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5641_ as2650.stack\[0\]\[9\] _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7921__A1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8360_ _3682_ _3697_ _3698_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4735__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ as2650.stack\[1\]\[5\] _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7311_ _1100_ _2582_ _2729_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4523_ _4102_ _4103_ _4104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8291_ _3635_ _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8477__A2 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7242_ _2661_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _3997_ _4034_ _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8709__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8229__A2 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _2586_ _2591_ _2593_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4385_ _3965_ _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6124_ _1054_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _1538_ _1426_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5006_ as2650.holding_reg\[5\] _0446_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_73_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4671__B1 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8401__A2 _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6412__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5215__A2 _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6957_ _1343_ _1305_ _2387_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5766__A3 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ _1375_ _1397_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6888_ _2321_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8627_ _0104_ clknet_3_0_0_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5839_ _1357_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7912__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4702__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__B1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8558_ _0035_ clknet_leaf_44_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6191__A3 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7509_ _2864_ _2886_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8489_ _2147_ _1370_ _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8468__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7140__A2 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7691__A3 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__I _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7979__A1 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5454__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__B1 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8156__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__A2 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7195__I _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7903__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5390__A1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8459__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5390__B2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5517__I0 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7131__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6890__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4496__A3 _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5445__A2 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6642__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7860_ _3248_ _3249_ _3250_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7198__A2 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8395__A1 _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6811_ _1288_ _2183_ _1371_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7791_ _3103_ _0643_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6945__A2 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6742_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4956__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8147__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6673_ _2132_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5618__I _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8412_ _0452_ _0455_ _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5624_ as2650.pc\[13\] _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4803__S1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8343_ _3683_ _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8531__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5381__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5555_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4506_ _3843_ as2650.ins_reg\[1\] _4087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8274_ _3616_ _3617_ _3618_ _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5486_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _2642_ _2644_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4437_ _4017_ _4011_ _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8681__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7156_ _2520_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4368_ _3864_ _3948_ _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6893__B _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6107_ _1314_ _3897_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7087_ _2220_ _2284_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4299_ as2650.cycle\[1\] _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6633__A1 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _0904_ _1517_ _0396_ _1554_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8386__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7989_ _3342_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6936__A2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4947__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5528__I _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7361__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5972__B _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__B2 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5911__A3 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7649__B1 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8310__A1 _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5124__A1 _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6872__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6624__A1 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A2 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8377__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8129__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7139__B _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__B _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5438__I _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__I _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5902__A3 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5340_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5271_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7010_ _1313_ _2170_ as2650.cycle\[2\] _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5666__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4469__A3 _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4874__B1 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6615__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7958__A4 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4517__I as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6091__A2 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7912_ _1133_ _1017_ _1264_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8368__A1 _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7843_ _1089_ _3239_ _3240_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5549__S _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4986_ _4160_ _0560_ _0585_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7774_ _1101_ _3100_ _3177_ _3129_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7591__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6725_ _2175_ _2176_ _1290_ _2177_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__I _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6656_ _2118_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _1155_ _1175_ _1176_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5354__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _0962_ _0865_ _2053_ _2033_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8326_ _3040_ _3667_ _3668_ _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _1077_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5106__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8257_ _2943_ _3602_ _3563_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5469_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5657__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7208_ _2621_ _2623_ _2627_ _2628_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_120_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8188_ _1547_ _0822_ _3535_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_115_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _2557_ _2559_ _2560_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6907__I _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8327__C _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5409__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6606__A1 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7231__C _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_55_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_100_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8577__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7031__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5593__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7334__A2 _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5896__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6089__I _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__A2 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8047__B1 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4320__A2 _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7270__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5820__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7022__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ _0341_ _0440_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7573__A2 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4771_ _0371_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ _1968_ _1974_ _1989_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7490_ _2903_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7325__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6441_ _4099_ _0528_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5336__A1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8479__I _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6501__B _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5887__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _1853_ _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8111_ _3441_ _3443_ _3447_ _3461_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7089__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5323_ _0881_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6836__A1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5639__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8042_ _0307_ _0331_ _3394_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_115_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5254_ _3886_ _3996_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7332__B _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6727__I _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ as2650.r0\[5\] _0367_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4862__A3 _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7261__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5811__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7826_ _2486_ _0803_ _2474_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5575__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _4000_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7757_ _0318_ _2214_ _1379_ _4223_ _3098_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_138_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ _2158_ _2161_ _2162_ _1359_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7688_ _1374_ _1412_ _2080_ _2229_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__6119__A3 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8513__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8513__B2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6639_ _2101_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5327__B2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5878__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4710__I _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__I1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8309_ _2367_ _2464_ _3648_ _3652_ _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4550__A2 _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4302__A2 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5541__I as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6055__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5802__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8504__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5318__A1 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5716__I _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5869__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4541__A2 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6818__A1 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5451__I _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7243__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6990_ _2418_ _2379_ _2419_ _2413_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7794__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5941_ _0290_ _4197_ _4053_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_59_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5872_ _3941_ _1319_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8660_ _0137_ clknet_leaf_71_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _4115_ _0416_ _0423_ _4118_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7611_ _2858_ _2996_ _3021_ _2682_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8591_ _0068_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__A3 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7542_ as2650.addr_buff\[1\] _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4754_ _4015_ _0346_ _0348_ _0350_ _0355_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8430__C _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7473_ _0713_ _0629_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4685_ as2650.r123\[1\]\[1\] _4253_ _0287_ _4155_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6424_ _0511_ _1658_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8510__A4 _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6355_ _0409_ _0741_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7841__I _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6809__A1 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5306_ _0897_ as2650.stack\[1\]\[8\] as2650.stack\[0\]\[8\] _0901_ _0902_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6286_ _1656_ _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_115_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8274__A3 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8025_ _3330_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5237_ _0677_ _0688_ _0695_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5361__I as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4296__A1 as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _0729_ _0760_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7234__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _0609_ _0694_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7785__A2 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6192__I _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7809_ _2486_ _0709_ _3209_ _3050_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8789_ _0266_ clknet_leaf_16_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8615__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4440__I _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4523__A2 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8765__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7751__I _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5271__I _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__A1 _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7700__B _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7776__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7926__I _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6051__B _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4470_ _3864_ _4050_ _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5011__I0 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7700__A2 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5711__A1 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6140_ _0840_ _1620_ _1629_ _1346_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6277__I _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6071_ _1103_ _1576_ _1583_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6806__A4 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4278__A1 _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _3923_ _0619_ _0620_ _0316_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__A2 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7610__B _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4953__C _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7767__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _2154_ _2398_ _2400_ _2403_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8712_ _0189_ clknet_leaf_30_wb_clk_i as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5924_ _0592_ _1441_ _0679_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__A1 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8643_ _0120_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5855_ _1372_ _1292_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8192__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _4101_ _0406_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8574_ _0051_ clknet_leaf_46_wb_clk_i as2650.stack\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8160__C _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5786_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7525_ _2937_ _2578_ _2938_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8788__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5950__A1 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4753__A2 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4737_ as2650.holding_reg\[2\] _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7456_ _2716_ as2650.stack\[1\]\[7\] as2650.stack\[0\]\[7\] _2758_ _2871_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4668_ _4067_ _4120_ _4247_ _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5389__S0 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8495__A3 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ _1846_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4505__A2 _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4599_ _4022_ _4178_ _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7387_ _2780_ _2782_ _2803_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_116_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6338_ as2650.r123_2\[2\]\[2\] _1717_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7504__C _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6258__A2 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6269_ _1722_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4269__A1 as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8008_ _3348_ _3356_ _3361_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7207__A1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6915__I _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7207__B2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__S _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7758__A2 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4441__A1 _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8183__A2 _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7930__A2 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5941__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5544__I1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5215__B _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7446__A1 _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7997__A2 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6825__I _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5472__A3 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6421__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8174__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6185__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _1065_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7921__A2 _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5571_ _1137_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4735__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _3856_ _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7310_ _2682_ _2728_ _2579_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _2854_ _2978_ _3503_ _3634_ _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7685__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7241_ _1364_ _1057_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4453_ _3918_ _4033_ _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7172_ _2592_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4384_ as2650.ins_reg\[5\] as2650.ins_reg\[6\] as2650.ins_reg\[7\] _3965_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7437__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ _3849_ _1620_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _1465_ _1525_ _1529_ _1505_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_85_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _0446_ _0538_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__A1 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__B2 _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__A2 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _3925_ _1282_ _2386_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5907_ _1403_ _1407_ _1419_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_34_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6887_ _2250_ _2324_ _2328_ _2092_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8165__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8626_ _0103_ clknet_leaf_1_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5838_ _4128_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8557_ _0034_ clknet_leaf_44_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5769_ _1287_ _4206_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7508_ as2650.pc\[8\] _2863_ _2886_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8488_ _3189_ _2360_ _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7439_ _2588_ _2842_ _2849_ _2853_ _2854_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5814__I _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7979__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8803__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6645__I as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6651__A2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__A1 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__A1 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__B2 _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6167__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7903__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5914__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7667__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5517__I1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7419__A1 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6890__A2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8092__A1 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5445__A3 _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6642__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8395__A2 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6810_ _1381_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7790_ _1109_ _3130_ _3192_ _3129_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6741_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8147__A2 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6672_ _2130_ _2131_ _2119_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8411_ _0486_ _0487_ _0510_ _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5623_ _1163_ _1189_ _1190_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8342_ _3683_ _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5554_ _1133_ _1064_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7658__A1 as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4505_ _4084_ _4085_ _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_8273_ _3570_ _3572_ _2322_ _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5485_ _1013_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7224_ _2643_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4436_ _4016_ as2650.carry _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6330__A1 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7155_ _2523_ _2571_ _2576_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4367_ _3940_ _3946_ _3947_ _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4892__A1 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6106_ _1315_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8083__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7086_ _1336_ _3961_ _2086_ _2250_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4298_ _3878_ _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7070__B _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6633__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7830__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6037_ as2650.psu\[3\] _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8386__A2 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7988_ _3315_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6939_ _0824_ _2364_ _2371_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8609_ _0086_ clknet_3_6_0_wb_clk_i as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__A1 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7649__B2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8310__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5124__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6872__A2 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6624__A2 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7821__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7821__B2 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4635__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8129__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4623__I _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6043__C _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6560__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8301__A2 _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5270_ _4131_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4874__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8065__A1 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6615__A2 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7812__A1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4626__A1 _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__C _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7911_ _3262_ _1252_ _3281_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8368__A2 _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6379__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7842_ as2650.stack\[6\]\[1\] _1602_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7576__B1 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7773_ _3101_ _3169_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4985_ as2650.r123\[1\]\[4\] _4253_ _0584_ _4154_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6724_ _1408_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7049__C _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6655_ _2088_ _2100_ _2106_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_118_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5606_ as2650.stack\[2\]\[10\] _1170_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6551__A1 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _2039_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8325_ _2180_ _1316_ _2615_ _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8256_ _2942_ _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6303__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5468_ _1052_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7207_ _0903_ as2650.stack\[3\]\[1\] as2650.stack\[2\]\[1\] _0906_ _2536_ _2628_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__6854__A2 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4419_ _3999_ _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8187_ _3512_ _3515_ _3534_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5399_ _0978_ _0934_ _0989_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7138_ _4065_ _2551_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6606__A2 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4708__I _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7803__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _2397_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6790__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5274__I _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8295__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8047__A1 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8047__B2 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4320__A3 _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__I _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4608__A1 _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7270__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5281__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6833__I _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6781__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _0289_ _4196_ _4156_ _4257_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_33_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8671__CLK clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6440_ _1917_ _1922_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6371_ _1776_ _1854_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8110_ _3453_ _3460_ _3321_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8286__A1 _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7089__A2 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5322_ _0866_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6836__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8041_ _3358_ _3392_ _3393_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5253_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7332__C _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5184_ _0746_ _0750_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__I _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7261__A2 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5272__A1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8210__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7013__A2 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7825_ _3133_ _0822_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5024__A1 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4263__I _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7756_ _1519_ _1501_ _2155_ _3160_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_40_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4968_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5575__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6707_ net24 _2158_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7687_ _2097_ _1039_ _2528_ _2234_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_123_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4899_ _0494_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8513__A2 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _2089_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6569_ _2038_ _1653_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8308_ _2493_ _3650_ _3651_ _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8277__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8239_ _2587_ _2914_ _3585_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6918__I _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8544__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5978__B _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8354__B _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A1 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7749__I as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__S0 _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5802__A3 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7004__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8201__A1 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5269__I _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6763__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5566__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8504__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5318__A2 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6818__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6828__I _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4348__I _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7243__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8440__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5940_ _0805_ _0799_ _1455_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_92_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5871_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5006__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7610_ _3019_ _3020_ _2273_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4822_ _4039_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6754__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8590_ _0067_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7541_ _2834_ _2946_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5021__A4 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4753_ _0351_ _0353_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7472_ _1129_ _2886_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4684_ _0286_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6423_ _0557_ _1759_ _1903_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8259__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6354_ _1747_ _1838_ _1795_ _1796_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__I _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6809__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6285_ _4195_ _1758_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8024_ _2145_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7062__C _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5236_ _0829_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _0734_ _0759_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7234__A2 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8431__A1 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5098_ _0433_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5245__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5796__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6993__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7808_ _2323_ _0706_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8788_ _0265_ clknet_leaf_15_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7739_ _3123_ _0392_ _3144_ _1471_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7170__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7473__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6984__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6736__A1 _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5539__A2 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5727__I _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8103__I _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4631__I _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8489__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7147__C _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5711__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ as2650.stack\[5\]\[3\] _1580_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ _0326_ _0313_ _0380_ _0493_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_113_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _2109_ _2269_ _2402_ _2142_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6975__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6975__B2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8711_ _0188_ clknet_leaf_30_wb_clk_i as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5923_ _0489_ _0491_ _0503_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8642_ _0119_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5854_ _0443_ _4133_ _0530_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4805_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _0298_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8573_ _0050_ clknet_leaf_45_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5785_ _1296_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7524_ _2166_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _0334_ _0337_ _4161_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5950__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7455_ _2757_ _2868_ _2869_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4667_ _3975_ as2650.idx_ctrl\[0\] _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ _1834_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7386_ _2548_ _2792_ _2802_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4598_ _4175_ _4177_ _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6337_ _1808_ _1821_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6268_ _1725_ _1754_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4269__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8007_ _3357_ _3359_ _3360_ _1708_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7801__B _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5219_ _4099_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6199_ _3938_ _1664_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5218__A1 _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7299__I _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7758__A3 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A2 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7766__I0 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7391__A1 _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4451__I _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5941__A2 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5154__B1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7446__A2 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5457__A1 _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7997__A3 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6957__A1 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4432__A2 _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7158__B _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6185__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7382__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4361__I _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5570_ _1112_ _1144_ _1145_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4521_ _4101_ _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7134__A1 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7240_ _2656_ _2658_ _2102_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7685__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4452_ _4009_ _4032_ _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5696__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _2391_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4383_ _3933_ _3963_ _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _1622_ _1337_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7437__A2 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6053_ _1497_ _1569_ _1469_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8605__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5004_ _4163_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6948__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6955_ _1058_ _1479_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8755__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5620__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5906_ _4204_ _1421_ _1423_ _1382_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_74_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6886_ _2325_ _2327_ _1434_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8625_ _0102_ clknet_leaf_35_wb_clk_i as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5837_ _1344_ _1355_ _1341_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7912__A3 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8556_ _0033_ clknet_leaf_44_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5923__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5768_ _3942_ _3914_ _3866_ _0354_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7507_ _2122_ _2920_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _4211_ _0303_ _0320_ _4208_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_136_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8487_ _3154_ _3809_ _3811_ _3813_ _2372_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7582__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7125__A1 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5699_ _1237_ _1230_ _1238_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7438_ _2306_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7515__C _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7369_ _0903_ as2650.stack\[3\]\[5\] as2650.stack\[2\]\[5\] _2540_ _2536_ _2786_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5830__I _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6100__A2 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6651__A3 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6939__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5611__A1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A2 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5277__I as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7492__I _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5127__B1 _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7667__A2 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5226__B _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4350__A1 _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8628__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8092__A2 _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5740__I _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8778__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8272__B _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6740_ _3991_ _1324_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6671_ as2650.addr_buff\[3\] _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8410_ _0605_ _0610_ _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5622_ as2650.stack\[2\]\[12\] _1170_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8341_ _3937_ _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5553_ _0884_ _1010_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4504_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _3854_ _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8272_ _3576_ _3578_ _1707_ _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5484_ _4055_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7223_ as2650.pc\[2\] net7 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4435_ as2650.psl\[3\] _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6330__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4341__A1 as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7154_ _2524_ _2575_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4366_ as2650.cycle\[1\] _3881_ _3878_ _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_116_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6105_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4892__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7085_ _2079_ _2476_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8083__A2 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ _3876_ _3877_ _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _1549_ _1551_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7830__A2 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4266__I _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8386__A3 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7987_ _2433_ _3341_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7594__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _2342_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _2305_ _1612_ _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8608_ _0085_ clknet_3_3_0_wb_clk_i as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7897__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8539_ _0016_ clknet_3_7_0_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5825__I _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7261__B _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6656__I _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8074__A2 _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__A2 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6388__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7337__A1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7888__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6560__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5470__I _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7812__A2 _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5823__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4626__A2 _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7910_ as2650.stack\[3\]\[14\] _1249_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7841_ _1593_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6379__A2 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7576__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7576__B2 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7772_ _0401_ _1625_ _1423_ _1900_ _3175_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4984_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ _1470_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6654_ _2107_ _2114_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7879__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6585_ _0961_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6551__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8324_ _2850_ _3663_ _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5536_ _1116_ _1085_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4562__A1 _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8255_ _3592_ _3594_ _3600_ _2461_ _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5467_ _4013_ _1053_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7206_ _0892_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4418_ as2650.r0\[0\] _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8186_ _1484_ _0706_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8177__B _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5398_ _0979_ _0936_ _0869_ _0988_ _0861_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7137_ _2102_ _2558_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4349_ _3890_ _3929_ _3897_ _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6067__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ _2402_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6019_ _4016_ _0395_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4925__S _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4724__I _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7100__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6790__A2 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A2 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5555__I _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A1 _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8295__A2 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8047__A2 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5290__I as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5223__C _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5281__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7558__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__I _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7730__A1 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4544__A1 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _1778_ _1803_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5321_ _0849_ _3991_ _4127_ _0916_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8286__A2 _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8040_ _1514_ _4244_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5252_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4809__I _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5183_ _0778_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6049__A1 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7797__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5272__A2 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7549__A1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8210__A2 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7824_ _1125_ _3130_ _3223_ _3224_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5024__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4967_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7755_ _3153_ _1900_ _3159_ _1501_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6706_ _2159_ _2160_ _2082_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4783__A1 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7686_ _3089_ _3092_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4898_ _0495_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6637_ _2093_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5375__I _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7721__A1 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6568_ _0864_ _2037_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8307_ _3005_ _3003_ _3625_ _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5519_ as2650.stack\[0\]\[3\] _1090_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6499_ _0825_ _1762_ _1979_ _1679_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8238_ _2881_ _3568_ _3503_ _2926_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8029__A2 _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8169_ _3350_ _3516_ _3517_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4697__S1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8201__A2 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A1 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7960__A1 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6763__A2 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8801__D _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5285__I _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7712__A1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6279__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A2 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4629__I _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7005__I _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7228__B1 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7779__A1 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8440__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5254__A2 _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5870_ _1385_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7400__B1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4821_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6754__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7951__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7540_ _2952_ _2922_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4752_ _3917_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6512__C _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7471_ _1123_ _2841_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4683_ _4258_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6506__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7703__A1 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _1760_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5128__C _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6353_ _0293_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7624__B _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5304_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6284_ _4249_ _1759_ _1769_ _1704_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_143_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8023_ _3343_ _3375_ _3376_ _3224_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5235_ _0678_ _0680_ _0685_ _0695_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4296__A3 as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6690__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5166_ _3992_ _0727_ _0763_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8431__A2 _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5097_ _0683_ _0635_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5245__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6993__A2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4274__I _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7807_ _3164_ _1976_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8190__B _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8787_ _0264_ clknet_leaf_15_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7942__A1 as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7585__I _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5999_ _0304_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7518__C _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7738_ _1478_ _4202_ _3142_ _3143_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7669_ _2636_ _3067_ _2682_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5038__C _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7170__A2 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6929__I _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7253__C _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6681__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8661__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6664__I _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6984__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8186__A1 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A2 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4912__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8489__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7444__B _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8110__A1 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5020_ _0326_ _0327_ _0380_ _0493_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_97_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6971_ _2401_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8710_ _0187_ clknet_leaf_36_wb_clk_i as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4986__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5922_ _0432_ _1439_ _0504_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8177__A1 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5853_ _3874_ _3932_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8641_ _0118_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4804_ _4105_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4738__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8572_ _0049_ clknet_leaf_45_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5784_ _1053_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7523_ _1157_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _0335_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8534__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7454_ as2650.stack\[6\]\[7\] _0907_ _2718_ as2650.stack\[7\]\[7\] _2869_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_120_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4666_ _4040_ _4245_ _4052_ _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6405_ _1878_ _1888_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7385_ _2701_ _2796_ _2801_ _2615_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5653__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4597_ _4009_ _4068_ _4025_ _4176_ _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8684__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7073__C _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6336_ _0363_ _1820_ _1695_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8101__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6267_ _1727_ _1753_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8006_ _1515_ _3357_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5218_ _4112_ _0805_ _0812_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _4111_ _1683_ _1684_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5149_ as2650.r0\[2\] _0565_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8404__A2 _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6415__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5218__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8168__A1 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6718__A2 _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5828__I _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7766__I1 _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7391__A2 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5941__A3 _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5154__A1 _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5154__B2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6654__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5457__A2 _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8159__A1 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8557__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__I _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6185__A3 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5393__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _4084_ _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8331__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7134__A2 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5145__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4451_ _4005_ _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7685__A3 _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6893__A1 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5696__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7170_ _2587_ _2588_ _2589_ _2590_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4382_ _3958_ _3962_ _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _1511_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _1531_ _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _0592_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__I _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6948__A2 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7070__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__A1 _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6954_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5905_ _1422_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6885_ _2326_ _2077_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8024__I _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8624_ _0101_ clknet_leaf_50_wb_clk_i as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5836_ _1345_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5767_ _1282_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8555_ _0032_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7506_ _2919_ _2890_ _2603_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4718_ _0308_ _4228_ _0319_ _4210_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8322__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8486_ _3738_ _3812_ _3671_ _0830_ _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5698_ as2650.stack\[2\]\[3\] _1235_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7125__A2 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7437_ _1639_ _2850_ _2852_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4649_ as2650.ins_reg\[5\] _3868_ as2650.ins_reg\[7\] _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _0892_ _2784_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6319_ _1719_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7299_ _0890_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6636__A1 _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8389__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5611__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5558__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7116__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5127__B2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6875__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6627__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7052__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4372__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6670_ _1520_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5366__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5366__B2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8340_ _3681_ _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5552_ _1105_ _1131_ _1132_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8304__A1 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4503_ _3857_ _3858_ _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8271_ _2122_ _2125_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5118__A1 _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5483_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4321__B _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7658__A3 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7222_ _2596_ _2640_ _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4434_ _4014_ _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7153_ _2573_ _2569_ _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4341__A2 _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4365_ _3941_ _3945_ _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6618__A1 _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6104_ _1377_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7084_ _2223_ _2231_ _2504_ _2505_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4296_ as2650.cycle\[7\] as2650.cycle\[6\] as2650.cycle\[5\] as2650.cycle\[4\] _3877_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_112_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8722__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4547__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6094__A2 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6035_ _0396_ _0398_ _0499_ _1508_ _1534_ _3847_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5841__A2 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7858__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7986_ _3307_ _3317_ _3340_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8182__C _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7594__A2 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7079__B _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6937_ _0808_ _2360_ _1526_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _2306_ _2307_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5357__A1 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8607_ _0084_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5819_ _3953_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7593__I _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ _3871_ _4070_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8538_ _0015_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5109__A1 _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8469_ _2448_ _0894_ _3796_ _3797_ _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6002__I _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6609__A1 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7282__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7034__A1 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5596__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4399__A2 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5288__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7337__A2 _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7717__B _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5899__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4920__I _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__B _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7008__I _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6848__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8745__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6076__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5823__A2 _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7840_ _1076_ _1600_ _3238_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__C _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7576__A2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7771_ _2130_ _1501_ _2155_ _3174_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4983_ _0578_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ _1316_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6653_ _1633_ _1625_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5604_ _0369_ _1156_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6584_ _1870_ _2028_ _2034_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8323_ _3592_ _3663_ _3665_ _2410_ _3149_ _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5535_ _1117_ _1084_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6839__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8254_ _3347_ _3599_ _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5466_ _3872_ _3943_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7205_ _2624_ as2650.stack\[1\]\[1\] as2650.stack\[0\]\[1\] _2625_ _2626_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4417_ _3997_ _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8185_ _2876_ _3532_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5397_ _0867_ _0985_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8177__C _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4348_ _3894_ _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7136_ net5 _4004_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4277__I as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7067_ _2434_ _2326_ _2479_ _2491_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_28_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4279_ _3859_ _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _0616_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6706__B _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7016__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7567__A2 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7969_ _3977_ _4124_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8618__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8212__I _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8768__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5750__A1 as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_33_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5571__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8507__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7730__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4544__A2 _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7961__I _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5320_ as2650.r123\[0\]\[0\] _0860_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8278__B _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6297__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _0521_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__I _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _4098_ _4002_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6049__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7246__A1 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7797__A2 _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7549__A2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7823_ _1358_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7754_ _1495_ _1472_ _3158_ _3121_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4966_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6705_ _1672_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7685_ _1083_ _3090_ _3091_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5656__I _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4897_ _0430_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6636_ _4130_ _2095_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4535__A2 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5732__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7871__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _1372_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8306_ _3649_ _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5518_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7804__C _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6498_ _1550_ _1670_ _1978_ _1667_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7485__A1 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8237_ _3565_ _3583_ _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5449_ _3892_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8168_ _1489_ _3354_ _3322_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7237__A1 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__B _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7119_ _2531_ as2650.stack\[5\]\[0\] as2650.stack\[4\]\[0\] _0898_ _2541_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5248__B1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8099_ _3448_ _3449_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7788__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__A3 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7960__A2 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4774__A2 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8590__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4526__A2 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7228__A1 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7730__B _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7228__B2 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7779__A2 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8440__A3 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4820_ _0419_ _0382_ _0385_ _0417_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7951__A2 _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _3981_ _0311_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5962__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7470_ _2548_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4682_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7703__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6421_ _0518_ _1810_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6352_ _0788_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7467__A1 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6283_ _4245_ _1690_ _1760_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8022_ net53 _3342_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5234_ _0426_ _0830_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7640__B _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4296__A4 as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5165_ as2650.r123\[1\]\[6\] _4151_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5096_ _4180_ _0681_ _0686_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5245__A3 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4453__A1 _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8471__B _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8195__A2 _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6770__I _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7806_ _1117_ _3100_ _3207_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8786_ _0263_ clknet_leaf_15_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7942__A2 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7737_ _1287_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4949_ _0543_ _3950_ _4210_ _0548_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7668_ _2471_ _3067_ _3074_ _3075_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6619_ _4048_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4508__A2 _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7599_ _2289_ _2712_ _3009_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7170__A3 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7534__C _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6010__I _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8806__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4995__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8186__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7933__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5944__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7697__A1 _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5172__A2 _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8110__A2 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4683__A1 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7621__A1 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__A2 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6970_ _1707_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _0343_ _1438_ _0437_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4986__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8177__A2 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8722__D _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8640_ _0117_ clknet_leaf_73_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5852_ _1286_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_34_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6188__A1 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7924__A2 _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ as2650.r123\[1\]\[4\] as2650.r123\[0\]\[4\] as2650.r123_2\[1\]\[4\] as2650.r123_2\[0\]\[4\]
+ _3844_ _0298_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8571_ _0048_ clknet_leaf_45_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4738__A2 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _1298_ _1300_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7522_ _2904_ _2918_ _2934_ _2935_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4734_ _4122_ _4222_ _0329_ _4120_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7688__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7453_ _0900_ as2650.stack\[5\]\[7\] as2650.stack\[4\]\[7\] _2758_ _2868_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4665_ _4244_ _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _1833_ _1887_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7384_ _1535_ _2384_ _2798_ _2800_ _2661_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4596_ _4008_ _4010_ _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6335_ _0337_ _1809_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8101__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6112__A1 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6266_ _1730_ _1752_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _1556_ _4245_ _3358_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7860__A1 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5217_ _4078_ _0813_ _4112_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6197_ _1661_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5148_ _0742_ _0743_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_111_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__A2 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7612__A1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5079_ as2650.holding_reg\[6\] _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6179__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5926__A1 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4729__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8769_ _0246_ clknet_leaf_31_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__C _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7679__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5844__I _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4901__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7300__B1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7280__B _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6654__A2 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5457__A3 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7603__A1 _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6624__B _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5090__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7439__C _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7906__A2 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5917__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6185__A4 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7119__B1 as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8331__A2 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6342__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4450_ _4015_ _4018_ _4030_ _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4381_ _3895_ _3961_ _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6893__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8095__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6120_ _1620_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6585__I _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _1532_ _1567_ _1526_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _0430_ _0495_ _0496_ _0491_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_67_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4408__A1 _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7070__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _2308_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5904_ _1413_ _4129_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6884_ _2075_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8623_ _0100_ clknet_leaf_49_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5908__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ as2650.psu\[5\] _1346_ _1349_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8554_ _0031_ clknet_leaf_57_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5384__A2 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8651__CLK clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6581__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _1008_ _1283_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7505_ _1546_ _4103_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7365__B _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _4227_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8485_ _1428_ _3737_ _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5697_ _1102_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ _2851_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4648_ _4227_ _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6333__A1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7367_ _2624_ as2650.stack\[1\]\[5\] as2650.stack\[0\]\[5\] _2531_ _2784_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4579_ _3992_ _4127_ _4152_ _4159_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_122_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8086__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ _1776_ _1778_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_104_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7298_ _2716_ as2650.stack\[5\]\[3\] as2650.stack\[4\]\[3\] _0895_ _2717_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6495__I _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8627__D _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _0745_ _0790_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8389__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5839__I _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8010__A1 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6572__A1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A2 _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6875__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A1 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8077__A1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6627__A2 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4918__I _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7824__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8524__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7052__A2 _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8674__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4810__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8001__A1 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7964__I _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__B1 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ _1185_ _1179_ _1187_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7185__B _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5551_ as2650.stack\[0\]\[7\] _1121_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8304__A2 _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _4081_ _4082_ _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8270_ _3559_ _3613_ _3615_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5118__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7658__A4 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7221_ as2650.pc\[1\] _1512_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4433_ _3982_ _4013_ _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7152_ _2469_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4364_ _3942_ _3944_ _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6618__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _1200_ _1600_ _1604_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7815__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4295_ as2650.cycle\[3\] as2650.cycle\[2\] _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7083_ _1388_ _1391_ _2184_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7204__I _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _1515_ _4185_ _0312_ _1517_ _0690_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4764__S _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8240__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8240__B2 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7985_ _1071_ _3318_ _3339_ _2174_ _3316_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5054__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _2364_ _2368_ _2369_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4801__A1 _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6867_ _2309_ _2263_ _1042_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8606_ _0083_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5818_ _1025_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6554__A1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6798_ _0635_ _0717_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8537_ _0014_ clknet_leaf_67_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5749_ _1234_ _1267_ _1273_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5109__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8468_ _0894_ _1295_ _2593_ _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7503__B1 _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7419_ _2834_ _2831_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8399_ _3730_ _1345_ _1478_ _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7806__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7114__I _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7282__A2 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__A1 as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6953__I _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8697__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7034__A2 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8231__A1 _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5045__A1 _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__I _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6793__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A1 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7742__B1 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8298__A1 _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6848__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7733__B _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6863__I _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5823__A3 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8222__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5479__I _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7770_ _3121_ _0614_ _3173_ _1411_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6784__A1 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _0579_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6721_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6812__B _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7694__I _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _1059_ _1029_ _1046_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5603_ _1172_ _1074_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6583_ as2650.r123_2\[0\]\[3\] _2045_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8289__A1 _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8322_ _3029_ _3664_ _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5534_ _0986_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_133_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6839__A2 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8253_ _3323_ _3596_ _3598_ _3103_ _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_106_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5465_ _3846_ _0521_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7204_ _0874_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8458__C _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4416_ _3995_ _3996_ _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8184_ _2877_ _3531_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _0986_ _0917_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4558__I _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7135_ _1511_ _4004_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4347_ _3889_ _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7066_ _2458_ _2487_ _2490_ _2374_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ _3857_ _3858_ _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7968_ _3322_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6919_ _2355_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7818__B _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7899_ _1248_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8516__A2 _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6527__A1 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7109__I _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6013__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5750__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4553__A3 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4468__I _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8452__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5266__A1 _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8204__A1 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__I _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5569__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6518__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8712__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7019__I _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5762__I as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5250_ _0466_ _0796_ _0846_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5181_ _0776_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8443__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7246__A2 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8725__D _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5009__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7822_ _3211_ _3222_ _3099_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6757__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7753_ _2038_ _3155_ _3157_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7638__B _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4965_ as2650.r123\[0\]\[4\] as2650.r123_2\[0\]\[4\] _0365_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6704_ _1464_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7684_ _2090_ _3966_ _4137_ _1046_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6509__B2 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__A2 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4896_ _0341_ _0440_ _0428_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6635_ _1707_ _2096_ _2097_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5032__I1 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7721__A3 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _1700_ _2027_ _2036_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5732__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8305_ _3005_ _3625_ _3003_ _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5517_ _1100_ _1101_ _1074_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6497_ _0718_ _1670_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8236_ _2410_ _3582_ _3168_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5448_ _3963_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5496__A1 _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4288__I _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8167_ _3512_ _3515_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5379_ _0924_ as2650.stack\[3\]\[12\] as2650.stack\[2\]\[12\] _0920_ _0971_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_120_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7237__A2 _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7118_ _0889_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8434__A1 _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8098_ _0393_ _0389_ _3386_ _3415_ _3416_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5248__B2 _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7049_ _1035_ _2103_ _2472_ _2475_ _2476_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_102_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5847__I _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8735__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7960__A3 _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7173__A1 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5723__A2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6920__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6678__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__B1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5582__I _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7228__A2 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5239__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4926__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8440__A4 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6739__A1 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7400__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _0339_ _3980_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5962__A2 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7164__A1 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ _4198_ _4158_ _4260_ _4153_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6420_ _1109_ _1663_ _1902_ _1860_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7703__A3 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _1832_ _1835_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5302_ _0872_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7467__A2 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6282_ _1086_ _1706_ _1767_ _1690_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8021_ _1082_ _3344_ _3373_ _3374_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5233_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8608__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5164_ _0465_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6978__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _0350_ _0689_ _0692_ _0349_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5650__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8758__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8854_ net47 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7805_ _3099_ _3206_ _2938_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8785_ _0262_ clknet_leaf_15_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7736_ _3140_ _3141_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4948_ _3949_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7667_ _0997_ _2675_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7155__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _0370_ _0371_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _3958_ _1039_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7815__C _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7598_ as2650.addr_buff\[3\] _2102_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4764__I0 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6549_ _0761_ _2016_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8219_ net35 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7831__B _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6969__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7630__A2 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__I _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7278__B _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A2 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7146__A1 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7697__A2 _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4380__A1 _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5880__A1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7621__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7967__I _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _1437_ _4175_ _0344_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ _0444_ _4133_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7385__A1 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6188__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4391__I _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4802_ _0397_ _4066_ _4074_ _0402_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_62_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8570_ _0047_ clknet_leaf_44_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5782_ as2650.psl\[7\] _0522_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5935__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7521_ _2522_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4733_ _4121_ _0324_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7137__A1 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7452_ _2863_ _2866_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7635__C _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4664_ _4067_ _4166_ _4243_ _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6403_ _1882_ _1886_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7383_ _2101_ _2799_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4595_ _4174_ _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6111__I _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6334_ _0331_ _1810_ _1697_ _1818_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6265_ _1735_ _1751_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6112__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8004_ _4063_ _4046_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5216_ as2650.psl\[3\] _4069_ _4017_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7860__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6196_ _1682_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8580__CLK clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5147_ _4079_ as2650.r0\[0\] _0525_ _0744_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7612__A2 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ _0628_ _0630_ _0632_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_56_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5623__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4426__A2 _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7376__A1 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6179__A2 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4515__B _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5926__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8768_ _0245_ clknet_leaf_32_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7826__B _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7719_ _3080_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8699_ _0176_ clknet_leaf_25_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7679__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7545__C _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6021__I as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7300__B2 as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7280__C _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7851__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5862__A1 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__A2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7367__A1 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7367__B2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7119__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7119__B2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4380_ _3905_ _3960_ _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6866__I _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _1334_ _1565_ _1566_ _1538_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7842__A2 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5853__A1 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A2 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _0592_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4386__I _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _2378_ _2382_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7070__A3 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5081__A2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5903_ _1420_ _1404_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6883_ _1463_ _2173_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6106__I _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8622_ _0099_ clknet_leaf_41_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5834_ _1346_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5010__I _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5908__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8553_ _0030_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ _0847_ _3973_ _0863_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5945__I _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4716_ _0312_ _0317_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7504_ _2905_ _2917_ _2527_ _2273_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8484_ _2159_ _3810_ _3809_ _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5696_ _1234_ _1230_ _1236_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7435_ _1315_ _2546_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _4226_ _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7530__A1 _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4344__A1 _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _2775_ _2780_ _2782_ _2470_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4578_ _4153_ _4155_ _4158_ _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4895__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6317_ _1779_ _1802_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8086__A2 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7297_ _0898_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ _1733_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6179_ _4072_ _1665_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6725__B _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7349__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8010__A2 _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_27_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8387__B _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6686__I _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6088__A1 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6635__B _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7588__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6260__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__A2 _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6012__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7185__C _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5550_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _3844_ _3858_ _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7512__A1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5118__A3 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4326__A1 as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7220_ as2650.pc\[1\] _1512_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4432_ _3869_ _4012_ _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6596__I _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7151_ _2572_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8068__A2 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4363_ _3914_ _3943_ _3944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6079__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ as2650.stack\[6\]\[14\] _1602_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7082_ _1362_ _1040_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7815__A2 _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _3874_ _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6033_ _0713_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7579__A1 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8240__A2 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7984_ _3320_ _3331_ _3338_ _1504_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6935_ _0683_ _2342_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4801__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6866_ _2308_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8605_ _0082_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5817_ _1031_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6797_ _0850_ _1303_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6554__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4565__A1 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8536_ _0013_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5748_ as2650.stack\[4\]\[2\] _1271_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ as2650.r123_2\[3\]\[5\] _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8467_ _3795_ _2345_ _2347_ _1344_ _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7503__B2 _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7418_ _4144_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8398_ _3729_ _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8059__A2 _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7349_ _2740_ _2756_ _2766_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7034__A3 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7130__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6793__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5585__I as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A2 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7742__A1 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7742__B2 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A1 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8298__A2 _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__I _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8641__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8222__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4981_ _0580_ _0577_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7981__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6784__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6720_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6812__C _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6651_ _1415_ _2112_ _2113_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_108_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6536__A2 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7733__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5495__I _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ as2650.pc\[10\] _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6582_ _2047_ _2050_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8321_ _3602_ _3025_ _3562_ _3027_ _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5533_ _1115_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8252_ _2955_ _3597_ _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6839__A3 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5464_ _3942_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7203_ _0872_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4415_ _3983_ _3915_ _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8183_ _2824_ _3510_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5395_ _0613_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7134_ _1070_ _2443_ _2553_ _2555_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4346_ as2650.addr_buff\[7\] _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7065_ _2109_ _2464_ _2489_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4277_ as2650.ins_reg\[1\] _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6016_ _1048_ _4014_ _1326_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A1 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7967_ _2112_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7972__A1 _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4786__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6918_ _2335_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7818__C _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7898_ _3248_ _3273_ _3274_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6849_ _1633_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6527__A2 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8519_ _3838_ _3840_ _1360_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8664__CLK clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8452__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5266__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__I _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8204__A2 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_42_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7963__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7715__A1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6204__I _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8140__A1 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ _0625_ _4255_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8443__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5257__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7651__B1 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4608__B _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6206__A1 _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ _0690_ _3137_ _3221_ _2267_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7954__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6757__A2 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4768__A1 _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4964_ _4213_ _0368_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7752_ _0369_ _3156_ _2674_ _0870_ _1477_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6703_ _2093_ _2145_ _2151_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__8537__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7683_ _1421_ _1422_ _1382_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4895_ as2650.holding_reg\[4\] _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7706__A1 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5980__A3 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6634_ _1413_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6565_ as2650.r123_2\[0\]\[0\] _2028_ _2030_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5953__I _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8304_ _3591_ _3641_ _3647_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5516_ _0962_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_121_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _0998_ _1662_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8131__A1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8235_ _3378_ _3568_ _3581_ _3347_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5447_ as2650.addr_buff\[7\] _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_47_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6693__A1 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5496__A2 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5378_ _0942_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8166_ _3478_ _3513_ _3514_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4329_ _3909_ _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7117_ _1020_ _2538_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8097_ _0394_ _0389_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7048_ _1547_ _1322_ _1611_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7642__B1 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8198__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__A2 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7945__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__I _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8370__A1 _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7173__A2 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6920__A2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__A1 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8122__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__B2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7476__A3 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6684__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7633__B1 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4998__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8189__A1 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6643__B _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5411__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _4259_ _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7164__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6350_ _1834_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8113__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4389__I _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6281_ _4202_ _1761_ _1766_ _1705_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8020_ _2174_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5232_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4525__I1 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5163_ _0729_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5094_ _0596_ _0690_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6978__A2 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__I _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5650__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8853_ net47 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7804_ _0540_ _3137_ _3195_ _3205_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_91_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8784_ _0261_ clknet_leaf_28_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5996_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7735_ _4260_ _2037_ _2629_ _3116_ _1494_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_40_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _0412_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7666_ _2696_ _3072_ _3073_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4878_ _0372_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6617_ _2074_ _2079_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5166__A1 _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7597_ _3004_ _3007_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4913__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4764__I1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6548_ _1949_ _2011_ _2021_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8104__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__I as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6479_ _1958_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6666__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8218_ _2493_ _3563_ _3564_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8149_ _2727_ _3498_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6969__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8702__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5641__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5858__I _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7918__A1 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7146__A2 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7294__B _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6689__I _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5157__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4904__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4380__A2 _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4507__I1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5880__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7606__B1 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7082__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7469__B _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _4102_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4801_ _3950_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5781_ _1299_ _0847_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5935__A3 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7520_ _0912_ _2529_ _2917_ _2933_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4732_ _4051_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8334__A1 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7451_ as2650.pc\[6\] _1114_ _2773_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4663_ _4067_ _4042_ _4242_ _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7688__A3 _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _1884_ _1885_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5699__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6896__A1 _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7382_ _2744_ _2746_ _2797_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4594_ as2650.holding_reg\[1\] _4090_ _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8098__B1 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6333_ _1687_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6648__A1 _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6264_ _1738_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_130_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6112__A3 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8003_ _3082_ _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5215_ _0808_ _4066_ _4211_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6195_ _1043_ _1493_ _1660_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_130_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _0740_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7073__A1 _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _3992_ _0649_ _0675_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5623__A2 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4582__I _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7376__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8767_ _0244_ clknet_leaf_32_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5979_ _1477_ _0804_ _1467_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7718_ _1622_ _1507_ _3122_ _3124_ _2694_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8698_ _0175_ clknet_leaf_25_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8325__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7128__A2 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7649_ _2931_ _3054_ _3057_ _2264_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7679__A3 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6887__A1 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7300__A2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__A2 _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6811__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5614__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5378__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6921__B _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8748__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5272__B _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ _0488_ _0491_ _0495_ _0505_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5853__A2 _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7055__A1 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6815__C _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6802__A1 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6802__B2 _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6951_ _2288_ _2379_ _2381_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__I _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5902_ _4021_ _1386_ _4164_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6882_ _2323_ _2081_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8621_ _0098_ clknet_leaf_41_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5833_ _4082_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_90_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8552_ _0029_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8307__A1 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _0461_ _4133_ _0523_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7503_ _2906_ _2904_ _2914_ _2915_ _2916_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4715_ _4092_ _4232_ _0314_ _0316_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4592__A2 _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8483_ _3730_ _2351_ _2350_ _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5695_ as2650.stack\[2\]\[2\] _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6869__A1 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7434_ _2551_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4646_ _3864_ _4145_ _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7530__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4344__A2 _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _4157_ _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7365_ _2781_ _2774_ _1312_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5961__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6316_ _1781_ _1801_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7296_ _2549_ _2700_ _2714_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4577__I _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6097__A2 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6247_ as2650.r0\[7\] _4256_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6178_ _3883_ _1664_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _4250_ _0698_ _0726_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_85_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6725__C _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7837__B _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__C _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_67_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5871__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8387__C _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6088__A2 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4487__I _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5835__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5820__B _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6260__A2 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5111__I _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7747__B _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6012__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5771__A1 _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8570__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4500_ _4080_ _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5480_ as2650.pc\[0\] _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7512__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6877__I _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4431_ _3915_ _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7150_ _1383_ _2288_ _2379_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4362_ as2650.ins_reg\[4\] _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6079__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6101_ _1194_ _1600_ _1603_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7276__A1 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7081_ _2319_ _2502_ _2503_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4293_ _3873_ _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _1547_ _0825_ _0539_ _0617_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7501__I _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7983_ _2304_ _3335_ _3337_ _1071_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6934_ _1125_ _1506_ _2367_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6865_ _1034_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5956__I _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6003__A2 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8604_ _0081_ clknet_leaf_54_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4860__I _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1027_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6796_ _2221_ _2223_ _2228_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__6280__C _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8535_ _0012_ clknet_leaf_65_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5747_ _1232_ _1267_ _1272_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8466_ _1352_ _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5678_ _1224_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7503__A2 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4317__A2 _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7417_ _2694_ _2565_ _2832_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4629_ _4208_ _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8397_ _0852_ _1351_ _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7348_ _2526_ _2739_ _2765_ _2630_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ _2683_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5817__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6736__B _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6793__A3 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8593__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5866__I _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6190__C _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7742__A2 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A2 _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6697__I _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7258__A1 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4867__I0 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7430__A1 _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4980_ _0478_ _0480_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7981__A2 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6381__B _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5992__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5776__I _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4680__I _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _1038_ _2076_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7196__C _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7733__A2 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5601_ _1155_ _1169_ _1171_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5744__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _0949_ _2032_ _2049_ _2040_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8320_ net40 _3662_ _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5532_ _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8251_ _2121_ _3570_ _3572_ _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5463_ _3963_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7202_ as2650.stack\[6\]\[1\] _2535_ _1015_ _2622_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4414_ _3994_ _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8182_ _3343_ _3529_ _3530_ _2435_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5394_ _0918_ _0980_ _0982_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7133_ _1030_ _2554_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _3903_ _3910_ _3925_ _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5016__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7064_ _2326_ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4276_ as2650.ins_reg\[0\] _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4855__I _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _1482_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7421__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6224__A2 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7966_ _2077_ _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ _2354_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4786__A2 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7897_ as2650.stack\[3\]\[8\] _1260_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5686__I _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4590__I _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6848_ _2288_ _2290_ _2258_ _2219_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6779_ _2184_ _2222_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_104_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8518_ _2362_ _3833_ _3839_ _3840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7488__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8449_ _2391_ _3143_ _1293_ _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5346__S0 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8452__A3 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4765__I _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7660__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6980__I _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7412__A1 as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7963__A2 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7715__A2 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7479__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__I _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4675__I _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__A3 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7651__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7651__B2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4465__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4608__C _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6206__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7403__A1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7820_ _2593_ _2242_ _3220_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7403__B2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7954__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7751_ _0853_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4768__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _0561_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6702_ _1398_ _2153_ _2154_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7682_ _1417_ _3088_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4894_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7706__A2 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6633_ _1377_ _1040_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5032__I3 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6564_ _0865_ _0912_ _2033_ _1072_ _2034_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__7654__C _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8303_ _3321_ _3644_ _3646_ _3366_ _2465_ _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5515_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6495_ _0698_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8131__A2 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6130__I _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8234_ _3103_ _3574_ _3580_ _3323_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5446_ _1027_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6693__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ _2844_ _0646_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5377_ _0921_ as2650.stack\[1\]\[12\] as2650.stack\[0\]\[12\] _0943_ _0969_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_87_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7116_ as2650.stack\[6\]\[0\] _0906_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4328_ _3908_ _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8096_ _3378_ _3446_ _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8057__I _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7642__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7047_ _2474_ _2413_ _2103_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7642__B2 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7896__I _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7945__A2 _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7949_ _1244_ _3286_ _3305_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8370__A2 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8631__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A2 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8122__A2 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6684__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7633__A1 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7633__B2 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4447__A1 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7800__S _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7739__C _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__B1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7046__I _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8113__A2 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5300_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6280_ _0392_ _1762_ _1765_ _1679_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5231_ _0826_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4686__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5162_ _0734_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__A1 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5093_ _0683_ _0596_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4989__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8852_ net47 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7927__A2 _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7803_ _2177_ _3196_ _3204_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8783_ _0260_ clknet_leaf_29_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7734_ _1443_ _3111_ _3139_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4946_ _3923_ _0513_ _0544_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8654__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4610__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7665__B _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7665_ _2587_ _2768_ _3067_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4877_ _0474_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5964__I _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8352__A2 _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8340__I _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6616_ _1413_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7384__C _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5166__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7596_ _3005_ _3006_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6547_ as2650.r123_2\[1\]\[5\] _2015_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8104__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6478_ _4099_ _1197_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8496__B _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6666__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8217_ _2907_ _3561_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5429_ _0897_ _1013_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8148_ _1116_ _3495_ _3496_ _3497_ _2780_ _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8079_ _2698_ _2389_ _2376_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7379__B1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7918__A2 _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__C _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8040__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__B2 _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5874__I _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7294__C _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__A2 _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4904__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7854__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A1 _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7606__A1 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8527__CLK clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7606__B2 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7082__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6654__B _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7469__C _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8677__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4840__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7909__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8031__A1 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4800_ _0398_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5396__A2 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5780_ as2650.psl\[7\] _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4731_ _4119_ _0323_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8334__A2 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7450_ _2864_ _2772_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4662_ _3934_ _4041_ _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7688__A4 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6401_ _0626_ _0527_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6896__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7381_ _2744_ _2746_ _2797_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4593_ _4170_ _4172_ _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6332_ _0290_ _1662_ _1815_ _1816_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8098__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6263_ _1742_ _1749_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__A1 _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8002_ _3350_ _3353_ _3355_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5214_ _4066_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6194_ _0291_ _1668_ _1677_ _1680_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5145_ _0561_ _0526_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__A2 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ as2650.r123\[1\]\[5\] _4151_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5959__I _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7379__C _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6283__C _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8022__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6584__A1 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8766_ _0243_ clknet_leaf_32_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5978_ _4097_ _1456_ _4024_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7717_ _3123_ _0291_ _1471_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4929_ _3844_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8697_ _0174_ clknet_leaf_25_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5694__I _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8325__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7648_ _3055_ _3056_ _2547_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7579_ _2935_ _2988_ _2990_ _2633_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_125_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7836__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8261__A1 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5075__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8245__I _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6811__A2 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4822__A1 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8013__A1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8013__B2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6575__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7772__B1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7752__C _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7827__A1 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8252__A1 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5066__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6950_ _2170_ _1383_ _2380_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6802__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4813__A1 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5901_ _0603_ _1330_ _1408_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__8004__A1 _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6881_ _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7994__I _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8620_ _0097_ clknet_leaf_41_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6566__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8551_ _0028_ clknet_leaf_57_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _4135_ _0854_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8307__A2 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7502_ _2302_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4714_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8482_ _3723_ _3724_ _3808_ _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5694_ _1153_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6869__A2 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7433_ _2843_ _2846_ _2848_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4645_ _4224_ _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5019__I _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4424__S0 _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7364_ _2564_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4576_ _4156_ _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6315_ _1783_ _1800_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7818__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4858__I _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7295_ _2701_ _2706_ _2713_ _2616_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_89_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8491__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _0749_ _1731_ _1732_ _0782_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ _3951_ _3850_ _4082_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_112_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _0334_ _0706_ _0725_ _4161_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _0657_ _0527_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8749_ _0226_ clknet_leaf_35_wb_clk_i as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7809__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8482__A1 _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6983__I _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8234__A1 _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8234__B2 _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5048__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6548__A1 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5771__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _4008_ _4010_ _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4361_ _3911_ _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6100_ as2650.stack\[6\]\[13\] _1602_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7080_ as2650.psu\[7\] _2319_ _2168_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7276__A2 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4292_ _3872_ _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _1539_ _4069_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7028__A2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7982_ _3336_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6787__A1 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5302__I _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _1606_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ net25 _2083_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8603_ _0080_ clknet_leaf_32_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5815_ _0530_ _1328_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6003__A3 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6795_ _2091_ _2188_ _2230_ _2238_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6133__I _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8534_ _0011_ clknet_leaf_65_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ as2650.stack\[4\]\[1\] _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4565__A3 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8465_ _3786_ _3793_ _0939_ _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5677_ as2650.r123_2\[3\]\[4\] _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7416_ _1612_ _2831_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4628_ _3903_ _4207_ _3988_ _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6711__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8396_ _1346_ _3718_ _3727_ _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7347_ _2761_ _2764_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4559_ _3927_ _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7267__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8464__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7278_ _2573_ _2695_ _2696_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7899__I _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5921__B _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6229_ _1368_ _1715_ _1654_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6736__C _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6778__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5450__A1 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8738__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8670__D _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6950__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5753__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6702__A1 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7750__I0 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8455__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4867__I1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8207__A1 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4492__A2 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6769__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5441__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7718__B1 _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5992__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5600_ as2650.stack\[2\]\[9\] _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6580_ _0948_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5744__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5531_ as2650.pc\[5\] _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5792__I _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8250_ _2955_ _3595_ _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5462_ _1030_ _1042_ _1047_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7201_ as2650.stack\[5\]\[1\] as2650.stack\[4\]\[1\] _0883_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4413_ _3913_ _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8181_ net34 _3342_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5393_ _0910_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7132_ _1068_ _4064_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8446__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4344_ _3919_ _3924_ _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7063_ as2650.cycle\[5\] _2480_ _3959_ _2438_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_115_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ _3855_ _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6014_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6128__I _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7421__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7965_ _3319_ _2554_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6572__B _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5967__I _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4871__I _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8343__I _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6916_ _0339_ _2352_ _2353_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7896_ _1251_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _1336_ _3961_ _2289_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7185__A1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6778_ _4048_ _1288_ _1290_ _1393_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6932__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5735__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8499__B _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5729_ _1239_ _1258_ _1259_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8517_ _3795_ _2361_ _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8448_ _1367_ _3773_ _3777_ _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8379_ net21 _3704_ _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5207__I _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8437__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6999__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5346__S1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8452__A4 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8560__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7412__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7176__A1 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5726__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8202__B _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7479__A2 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_51_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8428__A1 _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7636__C1 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4465__A2 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4691__I _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7954__A3 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4962_ _0468_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7750_ _0905_ _3154_ _3111_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6701_ _1290_ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7681_ _4049_ _3977_ _2225_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4893_ _0405_ _0407_ _0411_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6632_ _1044_ _1057_ _2094_ _2081_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5178__B1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6914__A1 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ _2029_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6390__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8302_ net39 _3645_ _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5514_ as2650.pc\[3\] _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6494_ _1968_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8233_ _2121_ _3579_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5445_ _1031_ _1032_ _3960_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5027__I _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7670__C _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8164_ _0615_ _0646_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7890__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ as2650.stack\[7\]\[12\] as2650.stack\[4\]\[12\] as2650.stack\[5\]\[12\] as2650.stack\[6\]\[12\]
+ _0938_ _0939_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7115_ _2534_ as2650.stack\[3\]\[0\] as2650.stack\[2\]\[0\] _2535_ _2536_ _2537_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4327_ _3906_ _3907_ _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8095_ net32 _3445_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7242__I _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _2473_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7642__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5697__I _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5405__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5405__B2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7948_ as2650.stack\[7\]\[6\] _3283_ _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7879_ _3262_ _1578_ _3263_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5708__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7330__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7881__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4695__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7152__I _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7633__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5644__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4447__A2 _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6991__I _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7397__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4725__B _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5400__I as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__B2 _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7755__C _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6372__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4383__A1 _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7771__B _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7321__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ as2650.holding_reg\[7\] _4109_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7872__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4525__I3 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5883__A1 _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4686__A2 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ _0738_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7624__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5092_ _0682_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__C _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8851_ net46 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7388__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7802_ _2136_ _1507_ _3197_ _3203_ _2392_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_92_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8782_ _0259_ clknet_leaf_28_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5994_ net6 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5310__I _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4945_ _0315_ _0314_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7733_ _0896_ _3138_ _0854_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A2 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7664_ _2446_ _3069_ _3071_ _2424_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4876_ _0475_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6615_ _2075_ _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7595_ _2974_ _2977_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7560__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6546_ _0673_ _2016_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7681__B _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6477_ _1883_ _1958_ _1923_ _1924_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_133_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8216_ _3562_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5428_ _1015_ _1010_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7863__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6910__I1 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8147_ _2389_ _2105_ _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5359_ _0935_ _0936_ _0933_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_47_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8078_ _3410_ _3412_ _3429_ _3149_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5626__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7029_ _2325_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7379__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4545__B _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7379__B2 _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8040__A2 _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5220__I _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7551__A1 _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4365__A1 _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5890__I _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7303__B2 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7854__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4507__I3 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7606__A2 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8031__A2 _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6042__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6593__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7790__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4730_ _4040_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4902__C _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4661_ _4198_ _4199_ _4201_ _4240_ _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_6400_ _1879_ _1883_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4356__A1 _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7380_ _0615_ _0534_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4592_ _4171_ _4091_ _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6331_ _0291_ _1682_ _1661_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8098__A2 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6262_ _1745_ _1748_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7845__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__A2 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5856__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8001_ _1516_ _3354_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5213_ _4108_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6193_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5305__I _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5144_ _3999_ _0741_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5075_ _0465_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6564__C _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6281__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8621__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8765_ _0242_ clknet_leaf_34_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7781__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5975__I _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8771__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7716_ _1467_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4928_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8696_ _0173_ clknet_leaf_20_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8325__A3 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7647_ _1191_ _3037_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7533__A1 _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4859_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_138_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7578_ _2968_ _2989_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _2007_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8300__B _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6739__C _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7836__A2 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7049__B1 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8261__A2 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__A3 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6046__I _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4822__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8013__A2 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6575__A2 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7772__A1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7772__B2 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__A1 _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7827__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8644__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7340__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5066__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4813__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5900_ _1412_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8004__A2 _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6880_ _2110_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ _1325_ _4143_ _1326_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5795__I _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5762_ as2650.psu\[5\] _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8550_ _0027_ clknet_leaf_57_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8307__A3 _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7501_ _2566_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4713_ _3866_ _3965_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7515__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8481_ _3774_ _1285_ _3807_ _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5693_ _1096_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4644_ net6 _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7432_ _2600_ _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4424__S1 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7363_ _2731_ _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4575_ _4002_ _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6314_ _1786_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7294_ _2709_ _2711_ _2712_ _2661_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7818__A2 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6245_ _0774_ _0783_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8491__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__I _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4501__A1 _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6176_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8346__I _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5127_ _3865_ _3901_ _4115_ _0709_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8243__A2 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5058_ as2650.r0\[0\] _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__A2 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6006__A1 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7754__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4568__A1 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8748_ _0225_ clknet_leaf_35_wb_clk_i as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7506__A1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8679_ _0156_ clknet_leaf_74_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4740__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7809__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7285__A3 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8482__A2 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8256__I _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_76_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6245__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5048__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A2 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6379__C _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4731__A1 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _3916_ _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4291_ as2650.ins_reg\[3\] _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6030_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6484__A1 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A2 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7981_ _1333_ _2249_ _2303_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7984__B2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6932_ _0586_ _2364_ _2366_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6863_ _1611_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8602_ _0079_ clknet_leaf_34_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5814_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__A4 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6794_ _2231_ _2232_ _2234_ _2237_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_50_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8533_ _0010_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5745_ _1268_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4970__A1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8464_ _1628_ _3766_ _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5676_ _1223_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7415_ _2824_ _2830_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4627_ _4206_ _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8395_ _3723_ _3724_ _3726_ _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6711__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4722__A1 _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4558_ _3956_ _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7346_ _2757_ _2762_ _2763_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4489_ _3921_ _4069_ _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7277_ _2469_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7672__B1 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _1704_ _1671_ _1714_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ _1648_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6227__A1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7975__A1 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6778__A2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5450__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6702__A2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7750__I1 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4713__A1 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6994__I _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput40 net40 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8207__A2 _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__A1 _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5441__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7718__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8391__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4952__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5530_ _1105_ _1112_ _1113_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8143__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4689__I _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5461_ _1048_ _4014_ _4143_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4412_ _3979_ _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7200_ as2650.stack\[7\]\[1\] _0878_ _1019_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8180_ _2812_ _3344_ _3528_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5392_ _0905_ as2650.stack\[3\]\[13\] as2650.stack\[2\]\[13\] _0908_ _0983_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_113_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7131_ _4065_ _2551_ _1416_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4343_ _3920_ _3923_ _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8446__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6457__A1 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7062_ _4140_ _2486_ _2293_ _1349_ _2227_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_119_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4274_ _3854_ _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _1493_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__A1 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7957__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7964_ _2397_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _2341_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7895_ _3262_ _1269_ _3272_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _1332_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7185__A2 _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8382__A1 _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7684__B _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6777_ _2217_ _2220_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5983__I _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8516_ _3814_ _3837_ as2650.psu\[4\] _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5728_ as2650.stack\[3\]\[4\] _1254_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8447_ _3774_ _1339_ _3776_ _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_87_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ as2650.stack\[1\]\[10\] _1213_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6696__A1 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8378_ _3700_ _4110_ _3712_ _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7329_ _2744_ _2745_ _2743_ _2710_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7645__B1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6999__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8705__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__A1 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6620__A1 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8373__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7176__A2 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8125__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6687__A1 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8428__A2 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7636__C2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5662__A2 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7769__B _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6611__A1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ as2650.r0\[1\] _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6700_ _1387_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7680_ _1502_ _2235_ _3926_ _3086_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4892_ _4170_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8364__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6631_ _1029_ _1034_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5178__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5178__B2 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6914__A2 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6562_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8116__A1 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8301_ _3628_ _3629_ _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5513_ _1067_ _1097_ _1098_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6493_ _1969_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5308__I _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8232_ _3576_ _3578_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5444_ _3905_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6848__B _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5350__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8163_ _1487_ _0705_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5350__B2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ _0870_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7114_ _1020_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4326_ as2650.cycle\[1\] _3896_ _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8094_ _3444_ _3413_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5102__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7045_ _2152_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6850__A1 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6602__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5405__A2 as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7947_ _1242_ _3286_ _3304_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7878_ as2650.stack\[5\]\[14\] _1575_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7158__A2 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6829_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4916__A1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8107__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6669__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__A1 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6841__A1 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5644__A2 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4792__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7397__A2 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__A2 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5837__B _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4907__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4383__A2 _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5580__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7771__C _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5332__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__B1 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5883__A2 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5160_ _0731_ _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7085__A1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5091_ _0677_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5635__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5798__I _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8850_ net46 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7388__A2 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7801_ _3121_ _3202_ _1471_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8781_ _0258_ clknet_leaf_29_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5993_ _4064_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7732_ _3110_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4944_ _4222_ _0302_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8337__A1 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7663_ _2422_ _3070_ _2931_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ _0294_ _4214_ _4156_ _4256_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_60_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6899__A1 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6614_ _2076_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7594_ as2650.pc\[10\] _1487_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6545_ _1909_ _2011_ _2019_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _0627_ _1957_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6578__B _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8215_ _2907_ _3561_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5427_ _1014_ _0890_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8146_ _2436_ _3475_ _2794_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5358_ _0871_ _0948_ _0950_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_47_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7076__A1 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4309_ as2650.cycle\[6\] _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8077_ _3410_ _3428_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5289_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7028_ _2440_ _2456_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7379__A2 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6587__B1 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A2 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7000__A1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7551__A2 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4365__A2 _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7591__C _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8500__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7067__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6814__A1 _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4736__B _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8319__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8573__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4660_ _4199_ _4239_ _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4356__A2 _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5553__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ as2650.holding_reg\[1\] _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _0398_ _1676_ _1814_ _1761_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6261_ _1743_ _1746_ _1747_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_143_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6648__A4 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8000_ _3349_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5856__A2 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5212_ _4230_ _0634_ _0799_ _0701_ _4205_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1678_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7058__A1 as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5143_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _0651_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6281__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6417__I _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8764_ _0241_ clknet_leaf_34_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5976_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5241__B1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7781__A2 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7715_ _1531_ _4111_ _3119_ _3121_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4927_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8695_ _0172_ clknet_leaf_15_wb_clk_i as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7248__I _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7646_ as2650.pc\[13\] _3037_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4858_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7577_ _2775_ _2986_ _2696_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5991__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4789_ _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ _1655_ _2006_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ _0617_ _1812_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4400__I _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7049__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5940__B _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8129_ _0617_ _1940_ _3478_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_48_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7221__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7772__A2 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4586__A2 _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6062__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4338__A2 _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7288__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5761_ _1246_ _1275_ _1280_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7068__I _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7500_ _2907_ _2913_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4712_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8480_ _3080_ _1519_ _2355_ _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5692_ _1232_ _1230_ _1233_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7515__A2 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7431_ _2843_ _2846_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4643_ _4222_ _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _2776_ _2778_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4574_ _4154_ _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _1789_ _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7293_ _1520_ _2604_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6244_ _0408_ _0566_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _4039_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7451__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5057_ _0570_ _0573_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7687__B _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__I _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8400__B1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8362__I _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4823__C _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7754__A2 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4568__A2 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8747_ _0224_ clknet_leaf_50_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5765__A1 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5959_ _4207_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8678_ _0155_ clknet_leaf_1_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7506__A2 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__B _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7629_ _3037_ _3038_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6190__A1 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4740__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__S0 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__I _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6796__A3 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5205__B1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5205__C2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7745__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8170__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8458__B1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4731__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4290_ _3867_ _3870_ _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7681__A1 _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6484__A2 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8761__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7980_ _2616_ _2554_ _3332_ _3334_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_82_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6931_ _2364_ _2365_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6862_ _1562_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8601_ _0078_ clknet_leaf_34_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5813_ _3947_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6793_ _1363_ _2235_ _2236_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_50_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8532_ _0009_ clknet_leaf_69_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5744_ _1228_ _1267_ _1270_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8463_ _1359_ _3785_ _3792_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5675_ as2650.r123_2\[3\]\[3\] _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8161__A2 _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7414_ _2825_ _2826_ _2829_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6172__A1 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4626_ _3942_ _4205_ _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8394_ _2147_ _2386_ _2498_ _3725_ _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6711__A3 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7345_ as2650.stack\[6\]\[4\] _2668_ _2718_ as2650.stack\[7\]\[4\] _0880_ _2763_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4557_ _3952_ _3956_ _4137_ _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4722__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7276_ _2639_ _2685_ _2693_ _2694_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4488_ _4068_ _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7672__A1 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _1687_ _1684_ _1702_ _1703_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ as2650.r123\[3\]\[5\] _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7424__A1 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6227__A2 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _4044_ _0700_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6089_ _1593_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7975__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6778__A3 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A1 _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6950__A3 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7436__I _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_opt_2_1_wb_clk_i clknet_opt_2_0_wb_clk_i clknet_opt_2_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8152__A2 _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6702__A3 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8784__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput30 net30 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7663__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4795__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7171__I _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__A1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7415__A1 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6218__A2 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7718__A2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5729__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4952__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8143__A2 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5460_ _3888_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _3849_ _3991_ _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7790__B _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5901__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5391_ _0941_ _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7130_ as2650.addr_buff\[0\] _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4342_ _3922_ _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8446__A3 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6457__A2 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7654__A1 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7061_ _2485_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4273_ _3853_ _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7654__B2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _1457_ _1455_ _1526_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
.ends

